VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MEM2_136X32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2_136X32 0 0 ;
  SIZE 422.725 BY 184.395 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 130.095 12.66 130.755 ;
      LAYER Metal6 ;
        RECT 12 130.095 12.66 130.755 ;
      LAYER Metal3 ;
        RECT 12 130.095 12.66 130.755 ;
      LAYER Metal4 ;
        RECT 12 130.095 12.66 130.755 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 123.975 12.66 124.635 ;
      LAYER Metal6 ;
        RECT 12 123.975 12.66 124.635 ;
      LAYER Metal3 ;
        RECT 12 123.975 12.66 124.635 ;
      LAYER Metal4 ;
        RECT 12 123.975 12.66 124.635 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 114.755 12.66 115.415 ;
      LAYER Metal6 ;
        RECT 12 114.755 12.66 115.415 ;
      LAYER Metal3 ;
        RECT 12 114.755 12.66 115.415 ;
      LAYER Metal4 ;
        RECT 12 114.755 12.66 115.415 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 111.735 12.66 112.395 ;
      LAYER Metal6 ;
        RECT 12 111.735 12.66 112.395 ;
      LAYER Metal3 ;
        RECT 12 111.735 12.66 112.395 ;
      LAYER Metal4 ;
        RECT 12 111.735 12.66 112.395 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 108.635 12.66 109.295 ;
      LAYER Metal6 ;
        RECT 12 108.635 12.66 109.295 ;
      LAYER Metal3 ;
        RECT 12 108.635 12.66 109.295 ;
      LAYER Metal4 ;
        RECT 12 108.635 12.66 109.295 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 102.515 12.66 103.175 ;
      LAYER Metal6 ;
        RECT 12 102.515 12.66 103.175 ;
      LAYER Metal3 ;
        RECT 12 102.515 12.66 103.175 ;
      LAYER Metal4 ;
        RECT 12 102.515 12.66 103.175 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 99.495 12.66 100.155 ;
      LAYER Metal6 ;
        RECT 12 99.495 12.66 100.155 ;
      LAYER Metal3 ;
        RECT 12 99.495 12.66 100.155 ;
      LAYER Metal4 ;
        RECT 12 99.495 12.66 100.155 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 96.395 12.66 97.055 ;
      LAYER Metal6 ;
        RECT 12 96.395 12.66 97.055 ;
      LAYER Metal3 ;
        RECT 12 96.395 12.66 97.055 ;
      LAYER Metal4 ;
        RECT 12 96.395 12.66 97.055 ;
    END
  END A1[7]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 51.835 12.66 52.495 ;
      LAYER Metal6 ;
        RECT 12 51.835 12.66 52.495 ;
      LAYER Metal3 ;
        RECT 12 51.835 12.66 52.495 ;
      LAYER Metal4 ;
        RECT 12 51.835 12.66 52.495 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 57.955 12.66 58.615 ;
      LAYER Metal6 ;
        RECT 12 57.955 12.66 58.615 ;
      LAYER Metal3 ;
        RECT 12 57.955 12.66 58.615 ;
      LAYER Metal4 ;
        RECT 12 57.955 12.66 58.615 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 67.175 12.66 67.835 ;
      LAYER Metal6 ;
        RECT 12 67.175 12.66 67.835 ;
      LAYER Metal3 ;
        RECT 12 67.175 12.66 67.835 ;
      LAYER Metal4 ;
        RECT 12 67.175 12.66 67.835 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 70.195 12.66 70.855 ;
      LAYER Metal6 ;
        RECT 12 70.195 12.66 70.855 ;
      LAYER Metal3 ;
        RECT 12 70.195 12.66 70.855 ;
      LAYER Metal4 ;
        RECT 12 70.195 12.66 70.855 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 73.295 12.66 73.955 ;
      LAYER Metal6 ;
        RECT 12 73.295 12.66 73.955 ;
      LAYER Metal3 ;
        RECT 12 73.295 12.66 73.955 ;
      LAYER Metal4 ;
        RECT 12 73.295 12.66 73.955 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 79.415 12.66 80.075 ;
      LAYER Metal6 ;
        RECT 12 79.415 12.66 80.075 ;
      LAYER Metal3 ;
        RECT 12 79.415 12.66 80.075 ;
      LAYER Metal4 ;
        RECT 12 79.415 12.66 80.075 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 82.435 12.66 83.095 ;
      LAYER Metal6 ;
        RECT 12 82.435 12.66 83.095 ;
      LAYER Metal3 ;
        RECT 12 82.435 12.66 83.095 ;
      LAYER Metal4 ;
        RECT 12 82.435 12.66 83.095 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 85.535 12.66 86.195 ;
      LAYER Metal6 ;
        RECT 12 85.535 12.66 86.195 ;
      LAYER Metal3 ;
        RECT 12 85.535 12.66 86.195 ;
      LAYER Metal4 ;
        RECT 12 85.535 12.66 86.195 ;
    END
  END A2[7]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 202.485 12 203.145 12.66 ;
      LAYER Metal6 ;
        RECT 202.485 12 203.145 12.66 ;
      LAYER Metal3 ;
        RECT 202.485 12 203.145 12.66 ;
      LAYER Metal4 ;
        RECT 202.485 12 203.145 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal6 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal3 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal4 ;
        RECT 196.36 12 197.02 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 211.11 12 211.77 12.66 ;
      LAYER Metal6 ;
        RECT 211.11 12 211.77 12.66 ;
      LAYER Metal3 ;
        RECT 211.11 12 211.77 12.66 ;
      LAYER Metal4 ;
        RECT 211.11 12 211.77 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal6 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal3 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal4 ;
        RECT 187.735 12 188.395 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal6 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal3 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal4 ;
        RECT 15.86 12 16.52 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal6 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal3 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal4 ;
        RECT 122.26 12 122.92 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal6 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal3 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal4 ;
        RECT 142.4 12 143.06 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal6 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal3 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal4 ;
        RECT 143.54 12 144.2 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal6 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal3 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal4 ;
        RECT 163.68 12 164.34 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal6 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal3 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal4 ;
        RECT 164.82 12 165.48 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal6 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal3 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal4 ;
        RECT 184.96 12 185.62 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 213.885 12 214.545 12.66 ;
      LAYER Metal6 ;
        RECT 213.885 12 214.545 12.66 ;
      LAYER Metal3 ;
        RECT 213.885 12 214.545 12.66 ;
      LAYER Metal4 ;
        RECT 213.885 12 214.545 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.025 12 234.685 12.66 ;
      LAYER Metal6 ;
        RECT 234.025 12 234.685 12.66 ;
      LAYER Metal3 ;
        RECT 234.025 12 234.685 12.66 ;
      LAYER Metal4 ;
        RECT 234.025 12 234.685 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 235.165 12 235.825 12.66 ;
      LAYER Metal6 ;
        RECT 235.165 12 235.825 12.66 ;
      LAYER Metal3 ;
        RECT 235.165 12 235.825 12.66 ;
      LAYER Metal4 ;
        RECT 235.165 12 235.825 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 255.305 12 255.965 12.66 ;
      LAYER Metal6 ;
        RECT 255.305 12 255.965 12.66 ;
      LAYER Metal3 ;
        RECT 255.305 12 255.965 12.66 ;
      LAYER Metal4 ;
        RECT 255.305 12 255.965 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal6 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal3 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal4 ;
        RECT 36 12 36.66 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 256.445 12 257.105 12.66 ;
      LAYER Metal6 ;
        RECT 256.445 12 257.105 12.66 ;
      LAYER Metal3 ;
        RECT 256.445 12 257.105 12.66 ;
      LAYER Metal4 ;
        RECT 256.445 12 257.105 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 276.585 12 277.245 12.66 ;
      LAYER Metal6 ;
        RECT 276.585 12 277.245 12.66 ;
      LAYER Metal3 ;
        RECT 276.585 12 277.245 12.66 ;
      LAYER Metal4 ;
        RECT 276.585 12 277.245 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 277.725 12 278.385 12.66 ;
      LAYER Metal6 ;
        RECT 277.725 12 278.385 12.66 ;
      LAYER Metal3 ;
        RECT 277.725 12 278.385 12.66 ;
      LAYER Metal4 ;
        RECT 277.725 12 278.385 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 297.865 12 298.525 12.66 ;
      LAYER Metal6 ;
        RECT 297.865 12 298.525 12.66 ;
      LAYER Metal3 ;
        RECT 297.865 12 298.525 12.66 ;
      LAYER Metal4 ;
        RECT 297.865 12 298.525 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 299.005 12 299.665 12.66 ;
      LAYER Metal6 ;
        RECT 299.005 12 299.665 12.66 ;
      LAYER Metal3 ;
        RECT 299.005 12 299.665 12.66 ;
      LAYER Metal4 ;
        RECT 299.005 12 299.665 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 319.145 12 319.805 12.66 ;
      LAYER Metal6 ;
        RECT 319.145 12 319.805 12.66 ;
      LAYER Metal3 ;
        RECT 319.145 12 319.805 12.66 ;
      LAYER Metal4 ;
        RECT 319.145 12 319.805 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 320.285 12 320.945 12.66 ;
      LAYER Metal6 ;
        RECT 320.285 12 320.945 12.66 ;
      LAYER Metal3 ;
        RECT 320.285 12 320.945 12.66 ;
      LAYER Metal4 ;
        RECT 320.285 12 320.945 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 340.425 12 341.085 12.66 ;
      LAYER Metal6 ;
        RECT 340.425 12 341.085 12.66 ;
      LAYER Metal3 ;
        RECT 340.425 12 341.085 12.66 ;
      LAYER Metal4 ;
        RECT 340.425 12 341.085 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 341.565 12 342.225 12.66 ;
      LAYER Metal6 ;
        RECT 341.565 12 342.225 12.66 ;
      LAYER Metal3 ;
        RECT 341.565 12 342.225 12.66 ;
      LAYER Metal4 ;
        RECT 341.565 12 342.225 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 361.705 12 362.365 12.66 ;
      LAYER Metal6 ;
        RECT 361.705 12 362.365 12.66 ;
      LAYER Metal3 ;
        RECT 361.705 12 362.365 12.66 ;
      LAYER Metal4 ;
        RECT 361.705 12 362.365 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal6 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal3 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal4 ;
        RECT 37.14 12 37.8 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 362.845 12 363.505 12.66 ;
      LAYER Metal6 ;
        RECT 362.845 12 363.505 12.66 ;
      LAYER Metal3 ;
        RECT 362.845 12 363.505 12.66 ;
      LAYER Metal4 ;
        RECT 362.845 12 363.505 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 382.985 12 383.645 12.66 ;
      LAYER Metal6 ;
        RECT 382.985 12 383.645 12.66 ;
      LAYER Metal3 ;
        RECT 382.985 12 383.645 12.66 ;
      LAYER Metal4 ;
        RECT 382.985 12 383.645 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal6 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal3 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal4 ;
        RECT 57.28 12 57.94 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal6 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal3 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal4 ;
        RECT 58.42 12 59.08 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal6 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal3 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal4 ;
        RECT 78.56 12 79.22 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal6 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal3 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal4 ;
        RECT 79.7 12 80.36 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal6 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal3 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal4 ;
        RECT 99.84 12 100.5 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal6 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal3 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal4 ;
        RECT 100.98 12 101.64 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal6 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal3 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal4 ;
        RECT 121.12 12 121.78 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal6 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal3 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal4 ;
        RECT 25.36 12 26.02 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal6 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal3 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal4 ;
        RECT 131.76 12 132.42 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal6 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal3 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal4 ;
        RECT 132.9 12 133.56 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal6 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal3 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal4 ;
        RECT 153.04 12 153.7 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal6 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal3 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal4 ;
        RECT 154.18 12 154.84 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal6 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal3 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal4 ;
        RECT 174.32 12 174.98 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal6 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal3 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal4 ;
        RECT 175.46 12 176.12 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 223.385 12 224.045 12.66 ;
      LAYER Metal6 ;
        RECT 223.385 12 224.045 12.66 ;
      LAYER Metal3 ;
        RECT 223.385 12 224.045 12.66 ;
      LAYER Metal4 ;
        RECT 223.385 12 224.045 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 224.525 12 225.185 12.66 ;
      LAYER Metal6 ;
        RECT 224.525 12 225.185 12.66 ;
      LAYER Metal3 ;
        RECT 224.525 12 225.185 12.66 ;
      LAYER Metal4 ;
        RECT 224.525 12 225.185 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 244.665 12 245.325 12.66 ;
      LAYER Metal6 ;
        RECT 244.665 12 245.325 12.66 ;
      LAYER Metal3 ;
        RECT 244.665 12 245.325 12.66 ;
      LAYER Metal4 ;
        RECT 244.665 12 245.325 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 245.805 12 246.465 12.66 ;
      LAYER Metal6 ;
        RECT 245.805 12 246.465 12.66 ;
      LAYER Metal3 ;
        RECT 245.805 12 246.465 12.66 ;
      LAYER Metal4 ;
        RECT 245.805 12 246.465 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal6 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal3 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal4 ;
        RECT 26.5 12 27.16 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 265.945 12 266.605 12.66 ;
      LAYER Metal6 ;
        RECT 265.945 12 266.605 12.66 ;
      LAYER Metal3 ;
        RECT 265.945 12 266.605 12.66 ;
      LAYER Metal4 ;
        RECT 265.945 12 266.605 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 267.085 12 267.745 12.66 ;
      LAYER Metal6 ;
        RECT 267.085 12 267.745 12.66 ;
      LAYER Metal3 ;
        RECT 267.085 12 267.745 12.66 ;
      LAYER Metal4 ;
        RECT 267.085 12 267.745 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 287.225 12 287.885 12.66 ;
      LAYER Metal6 ;
        RECT 287.225 12 287.885 12.66 ;
      LAYER Metal3 ;
        RECT 287.225 12 287.885 12.66 ;
      LAYER Metal4 ;
        RECT 287.225 12 287.885 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 288.365 12 289.025 12.66 ;
      LAYER Metal6 ;
        RECT 288.365 12 289.025 12.66 ;
      LAYER Metal3 ;
        RECT 288.365 12 289.025 12.66 ;
      LAYER Metal4 ;
        RECT 288.365 12 289.025 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 308.505 12 309.165 12.66 ;
      LAYER Metal6 ;
        RECT 308.505 12 309.165 12.66 ;
      LAYER Metal3 ;
        RECT 308.505 12 309.165 12.66 ;
      LAYER Metal4 ;
        RECT 308.505 12 309.165 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 309.645 12 310.305 12.66 ;
      LAYER Metal6 ;
        RECT 309.645 12 310.305 12.66 ;
      LAYER Metal3 ;
        RECT 309.645 12 310.305 12.66 ;
      LAYER Metal4 ;
        RECT 309.645 12 310.305 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 329.785 12 330.445 12.66 ;
      LAYER Metal6 ;
        RECT 329.785 12 330.445 12.66 ;
      LAYER Metal3 ;
        RECT 329.785 12 330.445 12.66 ;
      LAYER Metal4 ;
        RECT 329.785 12 330.445 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 330.925 12 331.585 12.66 ;
      LAYER Metal6 ;
        RECT 330.925 12 331.585 12.66 ;
      LAYER Metal3 ;
        RECT 330.925 12 331.585 12.66 ;
      LAYER Metal4 ;
        RECT 330.925 12 331.585 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 351.065 12 351.725 12.66 ;
      LAYER Metal6 ;
        RECT 351.065 12 351.725 12.66 ;
      LAYER Metal3 ;
        RECT 351.065 12 351.725 12.66 ;
      LAYER Metal4 ;
        RECT 351.065 12 351.725 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 352.205 12 352.865 12.66 ;
      LAYER Metal6 ;
        RECT 352.205 12 352.865 12.66 ;
      LAYER Metal3 ;
        RECT 352.205 12 352.865 12.66 ;
      LAYER Metal4 ;
        RECT 352.205 12 352.865 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal6 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal3 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal4 ;
        RECT 46.64 12 47.3 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 372.345 12 373.005 12.66 ;
      LAYER Metal6 ;
        RECT 372.345 12 373.005 12.66 ;
      LAYER Metal3 ;
        RECT 372.345 12 373.005 12.66 ;
      LAYER Metal4 ;
        RECT 372.345 12 373.005 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 373.485 12 374.145 12.66 ;
      LAYER Metal6 ;
        RECT 373.485 12 374.145 12.66 ;
      LAYER Metal3 ;
        RECT 373.485 12 374.145 12.66 ;
      LAYER Metal4 ;
        RECT 373.485 12 374.145 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal6 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal3 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal4 ;
        RECT 47.78 12 48.44 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal6 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal3 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal4 ;
        RECT 67.92 12 68.58 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal6 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal3 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal4 ;
        RECT 69.06 12 69.72 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal6 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal3 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal4 ;
        RECT 89.2 12 89.86 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal6 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal3 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal4 ;
        RECT 90.34 12 91 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal6 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal3 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal4 ;
        RECT 110.48 12 111.14 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal6 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal3 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal4 ;
        RECT 111.62 12 112.28 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal6 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal3 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal4 ;
        RECT 18.28 12 18.94 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal6 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal3 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal4 ;
        RECT 125.56 12 126.22 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal6 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal3 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal4 ;
        RECT 139.1 12 139.76 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal6 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal3 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal4 ;
        RECT 146.84 12 147.5 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal6 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal3 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal4 ;
        RECT 160.38 12 161.04 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal6 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal3 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal4 ;
        RECT 168.12 12 168.78 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal6 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal3 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal4 ;
        RECT 181.66 12 182.32 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 217.185 12 217.845 12.66 ;
      LAYER Metal6 ;
        RECT 217.185 12 217.845 12.66 ;
      LAYER Metal3 ;
        RECT 217.185 12 217.845 12.66 ;
      LAYER Metal4 ;
        RECT 217.185 12 217.845 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 230.725 12 231.385 12.66 ;
      LAYER Metal6 ;
        RECT 230.725 12 231.385 12.66 ;
      LAYER Metal3 ;
        RECT 230.725 12 231.385 12.66 ;
      LAYER Metal4 ;
        RECT 230.725 12 231.385 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 238.465 12 239.125 12.66 ;
      LAYER Metal6 ;
        RECT 238.465 12 239.125 12.66 ;
      LAYER Metal3 ;
        RECT 238.465 12 239.125 12.66 ;
      LAYER Metal4 ;
        RECT 238.465 12 239.125 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 252.005 12 252.665 12.66 ;
      LAYER Metal6 ;
        RECT 252.005 12 252.665 12.66 ;
      LAYER Metal3 ;
        RECT 252.005 12 252.665 12.66 ;
      LAYER Metal4 ;
        RECT 252.005 12 252.665 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal6 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal3 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal4 ;
        RECT 32.7 12 33.36 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 259.745 12 260.405 12.66 ;
      LAYER Metal6 ;
        RECT 259.745 12 260.405 12.66 ;
      LAYER Metal3 ;
        RECT 259.745 12 260.405 12.66 ;
      LAYER Metal4 ;
        RECT 259.745 12 260.405 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 273.285 12 273.945 12.66 ;
      LAYER Metal6 ;
        RECT 273.285 12 273.945 12.66 ;
      LAYER Metal3 ;
        RECT 273.285 12 273.945 12.66 ;
      LAYER Metal4 ;
        RECT 273.285 12 273.945 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 281.025 12 281.685 12.66 ;
      LAYER Metal6 ;
        RECT 281.025 12 281.685 12.66 ;
      LAYER Metal3 ;
        RECT 281.025 12 281.685 12.66 ;
      LAYER Metal4 ;
        RECT 281.025 12 281.685 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 294.565 12 295.225 12.66 ;
      LAYER Metal6 ;
        RECT 294.565 12 295.225 12.66 ;
      LAYER Metal3 ;
        RECT 294.565 12 295.225 12.66 ;
      LAYER Metal4 ;
        RECT 294.565 12 295.225 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 302.305 12 302.965 12.66 ;
      LAYER Metal6 ;
        RECT 302.305 12 302.965 12.66 ;
      LAYER Metal3 ;
        RECT 302.305 12 302.965 12.66 ;
      LAYER Metal4 ;
        RECT 302.305 12 302.965 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 315.845 12 316.505 12.66 ;
      LAYER Metal6 ;
        RECT 315.845 12 316.505 12.66 ;
      LAYER Metal3 ;
        RECT 315.845 12 316.505 12.66 ;
      LAYER Metal4 ;
        RECT 315.845 12 316.505 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 323.585 12 324.245 12.66 ;
      LAYER Metal6 ;
        RECT 323.585 12 324.245 12.66 ;
      LAYER Metal3 ;
        RECT 323.585 12 324.245 12.66 ;
      LAYER Metal4 ;
        RECT 323.585 12 324.245 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 337.125 12 337.785 12.66 ;
      LAYER Metal6 ;
        RECT 337.125 12 337.785 12.66 ;
      LAYER Metal3 ;
        RECT 337.125 12 337.785 12.66 ;
      LAYER Metal4 ;
        RECT 337.125 12 337.785 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 344.865 12 345.525 12.66 ;
      LAYER Metal6 ;
        RECT 344.865 12 345.525 12.66 ;
      LAYER Metal3 ;
        RECT 344.865 12 345.525 12.66 ;
      LAYER Metal4 ;
        RECT 344.865 12 345.525 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 358.405 12 359.065 12.66 ;
      LAYER Metal6 ;
        RECT 358.405 12 359.065 12.66 ;
      LAYER Metal3 ;
        RECT 358.405 12 359.065 12.66 ;
      LAYER Metal4 ;
        RECT 358.405 12 359.065 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal6 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal3 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal4 ;
        RECT 40.44 12 41.1 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.145 12 366.805 12.66 ;
      LAYER Metal6 ;
        RECT 366.145 12 366.805 12.66 ;
      LAYER Metal3 ;
        RECT 366.145 12 366.805 12.66 ;
      LAYER Metal4 ;
        RECT 366.145 12 366.805 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 380.565 12 381.225 12.66 ;
      LAYER Metal6 ;
        RECT 380.565 12 381.225 12.66 ;
      LAYER Metal3 ;
        RECT 380.565 12 381.225 12.66 ;
      LAYER Metal4 ;
        RECT 380.565 12 381.225 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal6 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal3 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal4 ;
        RECT 53.98 12 54.64 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal6 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal3 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal4 ;
        RECT 61.72 12 62.38 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal6 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal3 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal4 ;
        RECT 75.26 12 75.92 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal6 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal3 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal4 ;
        RECT 83 12 83.66 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal6 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal3 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal4 ;
        RECT 96.54 12 97.2 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal6 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal3 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal4 ;
        RECT 104.28 12 104.94 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal6 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal3 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal4 ;
        RECT 117.82 12 118.48 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal6 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal3 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal4 ;
        RECT 22.06 12 22.72 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal6 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal3 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal4 ;
        RECT 128.46 12 129.12 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal6 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal3 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal4 ;
        RECT 136.2 12 136.86 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal6 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal3 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal4 ;
        RECT 149.74 12 150.4 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal6 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal3 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal4 ;
        RECT 157.48 12 158.14 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal6 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal3 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal4 ;
        RECT 171.02 12 171.68 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal6 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal3 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal4 ;
        RECT 178.76 12 179.42 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 220.085 12 220.745 12.66 ;
      LAYER Metal6 ;
        RECT 220.085 12 220.745 12.66 ;
      LAYER Metal3 ;
        RECT 220.085 12 220.745 12.66 ;
      LAYER Metal4 ;
        RECT 220.085 12 220.745 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 227.825 12 228.485 12.66 ;
      LAYER Metal6 ;
        RECT 227.825 12 228.485 12.66 ;
      LAYER Metal3 ;
        RECT 227.825 12 228.485 12.66 ;
      LAYER Metal4 ;
        RECT 227.825 12 228.485 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 241.365 12 242.025 12.66 ;
      LAYER Metal6 ;
        RECT 241.365 12 242.025 12.66 ;
      LAYER Metal3 ;
        RECT 241.365 12 242.025 12.66 ;
      LAYER Metal4 ;
        RECT 241.365 12 242.025 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 249.105 12 249.765 12.66 ;
      LAYER Metal6 ;
        RECT 249.105 12 249.765 12.66 ;
      LAYER Metal3 ;
        RECT 249.105 12 249.765 12.66 ;
      LAYER Metal4 ;
        RECT 249.105 12 249.765 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal6 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal3 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal4 ;
        RECT 29.8 12 30.46 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 262.645 12 263.305 12.66 ;
      LAYER Metal6 ;
        RECT 262.645 12 263.305 12.66 ;
      LAYER Metal3 ;
        RECT 262.645 12 263.305 12.66 ;
      LAYER Metal4 ;
        RECT 262.645 12 263.305 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 270.385 12 271.045 12.66 ;
      LAYER Metal6 ;
        RECT 270.385 12 271.045 12.66 ;
      LAYER Metal3 ;
        RECT 270.385 12 271.045 12.66 ;
      LAYER Metal4 ;
        RECT 270.385 12 271.045 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 283.925 12 284.585 12.66 ;
      LAYER Metal6 ;
        RECT 283.925 12 284.585 12.66 ;
      LAYER Metal3 ;
        RECT 283.925 12 284.585 12.66 ;
      LAYER Metal4 ;
        RECT 283.925 12 284.585 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.665 12 292.325 12.66 ;
      LAYER Metal6 ;
        RECT 291.665 12 292.325 12.66 ;
      LAYER Metal3 ;
        RECT 291.665 12 292.325 12.66 ;
      LAYER Metal4 ;
        RECT 291.665 12 292.325 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 305.205 12 305.865 12.66 ;
      LAYER Metal6 ;
        RECT 305.205 12 305.865 12.66 ;
      LAYER Metal3 ;
        RECT 305.205 12 305.865 12.66 ;
      LAYER Metal4 ;
        RECT 305.205 12 305.865 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 312.945 12 313.605 12.66 ;
      LAYER Metal6 ;
        RECT 312.945 12 313.605 12.66 ;
      LAYER Metal3 ;
        RECT 312.945 12 313.605 12.66 ;
      LAYER Metal4 ;
        RECT 312.945 12 313.605 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 326.485 12 327.145 12.66 ;
      LAYER Metal6 ;
        RECT 326.485 12 327.145 12.66 ;
      LAYER Metal3 ;
        RECT 326.485 12 327.145 12.66 ;
      LAYER Metal4 ;
        RECT 326.485 12 327.145 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 334.225 12 334.885 12.66 ;
      LAYER Metal6 ;
        RECT 334.225 12 334.885 12.66 ;
      LAYER Metal3 ;
        RECT 334.225 12 334.885 12.66 ;
      LAYER Metal4 ;
        RECT 334.225 12 334.885 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 347.765 12 348.425 12.66 ;
      LAYER Metal6 ;
        RECT 347.765 12 348.425 12.66 ;
      LAYER Metal3 ;
        RECT 347.765 12 348.425 12.66 ;
      LAYER Metal4 ;
        RECT 347.765 12 348.425 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 355.505 12 356.165 12.66 ;
      LAYER Metal6 ;
        RECT 355.505 12 356.165 12.66 ;
      LAYER Metal3 ;
        RECT 355.505 12 356.165 12.66 ;
      LAYER Metal4 ;
        RECT 355.505 12 356.165 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal6 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal3 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal4 ;
        RECT 43.34 12 44 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 369.045 12 369.705 12.66 ;
      LAYER Metal6 ;
        RECT 369.045 12 369.705 12.66 ;
      LAYER Metal3 ;
        RECT 369.045 12 369.705 12.66 ;
      LAYER Metal4 ;
        RECT 369.045 12 369.705 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.785 12 377.445 12.66 ;
      LAYER Metal6 ;
        RECT 376.785 12 377.445 12.66 ;
      LAYER Metal3 ;
        RECT 376.785 12 377.445 12.66 ;
      LAYER Metal4 ;
        RECT 376.785 12 377.445 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal6 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal3 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal4 ;
        RECT 51.08 12 51.74 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal6 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal3 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal4 ;
        RECT 64.62 12 65.28 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal6 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal3 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal4 ;
        RECT 72.36 12 73.02 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal6 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal3 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal4 ;
        RECT 85.9 12 86.56 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal6 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal3 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal4 ;
        RECT 93.64 12 94.3 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal6 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal3 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal4 ;
        RECT 107.18 12 107.84 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal6 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal3 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal4 ;
        RECT 114.92 12 115.58 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 204.885 12 205.545 12.66 ;
      LAYER Metal6 ;
        RECT 204.885 12 205.545 12.66 ;
      LAYER Metal3 ;
        RECT 204.885 12 205.545 12.66 ;
      LAYER Metal4 ;
        RECT 204.885 12 205.545 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal6 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal3 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal4 ;
        RECT 193.96 12 194.62 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 179.395 422.725 184.395 ;
        RECT 0 0 422.725 5 ;
      LAYER Metal2 ;
        RECT 417.725 0 422.725 184.395 ;
        RECT 0 0 5 184.395 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 173.795 417.125 178.795 ;
        RECT 5.6 5.6 417.125 10.6 ;
      LAYER Metal2 ;
        RECT 412.125 5.6 417.125 178.795 ;
        RECT 5.6 5.6 10.6 178.795 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 410.735 172.39 ;
    LAYER Metal2 ;
      RECT 12 12 410.735 172.39 ;
    LAYER Metal3 ;
      RECT 12 12 410.735 172.39 ;
    LAYER Metal4 ;
      RECT 12 12 410.735 172.39 ;
    LAYER Metal5 ;
      RECT 12 12 410.735 172.39 ;
    LAYER Metal6 ;
      RECT 12 12 410.735 172.39 ;
  END
END MEM2_136X32

END LIBRARY
