VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MEM2_512X32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2_512X32 0 0 ;
  SIZE 763.02 BY 207.2 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 147.55 12.66 148.21 ;
      LAYER Metal6 ;
        RECT 12 147.55 12.66 148.21 ;
      LAYER Metal3 ;
        RECT 12 147.55 12.66 148.21 ;
      LAYER Metal4 ;
        RECT 12 147.55 12.66 148.21 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 141.43 12.66 142.09 ;
      LAYER Metal6 ;
        RECT 12 141.43 12.66 142.09 ;
      LAYER Metal3 ;
        RECT 12 141.43 12.66 142.09 ;
      LAYER Metal4 ;
        RECT 12 141.43 12.66 142.09 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 138.33 12.66 138.99 ;
      LAYER Metal6 ;
        RECT 12 138.33 12.66 138.99 ;
      LAYER Metal3 ;
        RECT 12 138.33 12.66 138.99 ;
      LAYER Metal4 ;
        RECT 12 138.33 12.66 138.99 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 132.21 12.66 132.87 ;
      LAYER Metal6 ;
        RECT 12 132.21 12.66 132.87 ;
      LAYER Metal3 ;
        RECT 12 132.21 12.66 132.87 ;
      LAYER Metal4 ;
        RECT 12 132.21 12.66 132.87 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 129.19 12.66 129.85 ;
      LAYER Metal6 ;
        RECT 12 129.19 12.66 129.85 ;
      LAYER Metal3 ;
        RECT 12 129.19 12.66 129.85 ;
      LAYER Metal4 ;
        RECT 12 129.19 12.66 129.85 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 126.09 12.66 126.75 ;
      LAYER Metal6 ;
        RECT 12 126.09 12.66 126.75 ;
      LAYER Metal3 ;
        RECT 12 126.09 12.66 126.75 ;
      LAYER Metal4 ;
        RECT 12 126.09 12.66 126.75 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 119.97 12.66 120.63 ;
      LAYER Metal6 ;
        RECT 12 119.97 12.66 120.63 ;
      LAYER Metal3 ;
        RECT 12 119.97 12.66 120.63 ;
      LAYER Metal4 ;
        RECT 12 119.97 12.66 120.63 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 116.95 12.66 117.61 ;
      LAYER Metal6 ;
        RECT 12 116.95 12.66 117.61 ;
      LAYER Metal3 ;
        RECT 12 116.95 12.66 117.61 ;
      LAYER Metal4 ;
        RECT 12 116.95 12.66 117.61 ;
    END
  END A1[7]
  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 113.85 12.66 114.51 ;
      LAYER Metal6 ;
        RECT 12 113.85 12.66 114.51 ;
      LAYER Metal3 ;
        RECT 12 113.85 12.66 114.51 ;
      LAYER Metal4 ;
        RECT 12 113.85 12.66 114.51 ;
    END
  END A1[8]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 69.29 12.66 69.95 ;
      LAYER Metal6 ;
        RECT 12 69.29 12.66 69.95 ;
      LAYER Metal3 ;
        RECT 12 69.29 12.66 69.95 ;
      LAYER Metal4 ;
        RECT 12 69.29 12.66 69.95 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 75.41 12.66 76.07 ;
      LAYER Metal6 ;
        RECT 12 75.41 12.66 76.07 ;
      LAYER Metal3 ;
        RECT 12 75.41 12.66 76.07 ;
      LAYER Metal4 ;
        RECT 12 75.41 12.66 76.07 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 78.51 12.66 79.17 ;
      LAYER Metal6 ;
        RECT 12 78.51 12.66 79.17 ;
      LAYER Metal3 ;
        RECT 12 78.51 12.66 79.17 ;
      LAYER Metal4 ;
        RECT 12 78.51 12.66 79.17 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 84.63 12.66 85.29 ;
      LAYER Metal6 ;
        RECT 12 84.63 12.66 85.29 ;
      LAYER Metal3 ;
        RECT 12 84.63 12.66 85.29 ;
      LAYER Metal4 ;
        RECT 12 84.63 12.66 85.29 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 87.65 12.66 88.31 ;
      LAYER Metal6 ;
        RECT 12 87.65 12.66 88.31 ;
      LAYER Metal3 ;
        RECT 12 87.65 12.66 88.31 ;
      LAYER Metal4 ;
        RECT 12 87.65 12.66 88.31 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 90.75 12.66 91.41 ;
      LAYER Metal6 ;
        RECT 12 90.75 12.66 91.41 ;
      LAYER Metal3 ;
        RECT 12 90.75 12.66 91.41 ;
      LAYER Metal4 ;
        RECT 12 90.75 12.66 91.41 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 96.87 12.66 97.53 ;
      LAYER Metal6 ;
        RECT 12 96.87 12.66 97.53 ;
      LAYER Metal3 ;
        RECT 12 96.87 12.66 97.53 ;
      LAYER Metal4 ;
        RECT 12 96.87 12.66 97.53 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 99.89 12.66 100.55 ;
      LAYER Metal6 ;
        RECT 12 99.89 12.66 100.55 ;
      LAYER Metal3 ;
        RECT 12 99.89 12.66 100.55 ;
      LAYER Metal4 ;
        RECT 12 99.89 12.66 100.55 ;
    END
  END A2[7]
  PIN A2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 102.99 12.66 103.65 ;
      LAYER Metal6 ;
        RECT 12 102.99 12.66 103.65 ;
      LAYER Metal3 ;
        RECT 12 102.99 12.66 103.65 ;
      LAYER Metal4 ;
        RECT 12 102.99 12.66 103.65 ;
    END
  END A2[8]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 377.5 12.00 378.16 12.66 ;
      LAYER Metal6 ;
        RECT 377.5 12.00 378.16 12.66 ;
      LAYER Metal3 ;
        RECT 377.5 12.00 378.16 12.66 ;
      LAYER Metal4 ;
        RECT 377.5 12.00 378.16 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.6 12.00 367.26 12.66 ;
      LAYER Metal6 ;
        RECT 366.6 12.00 367.26 12.66 ;
      LAYER Metal3 ;
        RECT 366.6 12.00 367.26 12.66 ;
      LAYER Metal4 ;
        RECT 366.6 12.00 367.26 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 386.125 12.00 386.785 12.66 ;
      LAYER Metal6 ;
        RECT 386.125 12.00 386.785 12.66 ;
      LAYER Metal3 ;
        RECT 386.125 12.00 386.785 12.66 ;
      LAYER Metal4 ;
        RECT 386.125 12.00 386.785 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 357.975 12.00 358.635 12.66 ;
      LAYER Metal6 ;
        RECT 357.975 12.00 358.635 12.66 ;
      LAYER Metal3 ;
        RECT 357.975 12.00 358.635 12.66 ;
      LAYER Metal4 ;
        RECT 357.975 12.00 358.635 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 21.91 12.00 22.57 12.66 ;
      LAYER Metal6 ;
        RECT 21.91 12.00 22.57 12.66 ;
      LAYER Metal3 ;
        RECT 21.91 12.00 22.57 12.66 ;
      LAYER Metal4 ;
        RECT 21.91 12.00 22.57 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.71 12.00 235.37 12.66 ;
      LAYER Metal6 ;
        RECT 234.71 12.00 235.37 12.66 ;
      LAYER Metal3 ;
        RECT 234.71 12.00 235.37 12.66 ;
      LAYER Metal4 ;
        RECT 234.71 12.00 235.37 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.03 12.00 264.69 12.66 ;
      LAYER Metal6 ;
        RECT 264.03 12.00 264.69 12.66 ;
      LAYER Metal3 ;
        RECT 264.03 12.00 264.69 12.66 ;
      LAYER Metal4 ;
        RECT 264.03 12.00 264.69 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 277.27 12.00 277.93 12.66 ;
      LAYER Metal6 ;
        RECT 277.27 12.00 277.93 12.66 ;
      LAYER Metal3 ;
        RECT 277.27 12.00 277.93 12.66 ;
      LAYER Metal4 ;
        RECT 277.27 12.00 277.93 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.59 12.00 307.25 12.66 ;
      LAYER Metal6 ;
        RECT 306.59 12.00 307.25 12.66 ;
      LAYER Metal3 ;
        RECT 306.59 12.00 307.25 12.66 ;
      LAYER Metal4 ;
        RECT 306.59 12.00 307.25 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 319.83 12.00 320.49 12.66 ;
      LAYER Metal6 ;
        RECT 319.83 12.00 320.49 12.66 ;
      LAYER Metal3 ;
        RECT 319.83 12.00 320.49 12.66 ;
      LAYER Metal4 ;
        RECT 319.83 12.00 320.49 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.15 12.00 349.81 12.66 ;
      LAYER Metal6 ;
        RECT 349.15 12.00 349.81 12.66 ;
      LAYER Metal3 ;
        RECT 349.15 12.00 349.81 12.66 ;
      LAYER Metal4 ;
        RECT 349.15 12.00 349.81 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 394.95 12.00 395.61 12.66 ;
      LAYER Metal6 ;
        RECT 394.95 12.00 395.61 12.66 ;
      LAYER Metal3 ;
        RECT 394.95 12.00 395.61 12.66 ;
      LAYER Metal4 ;
        RECT 394.95 12.00 395.61 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 424.27 12.00 424.93 12.66 ;
      LAYER Metal6 ;
        RECT 424.27 12.00 424.93 12.66 ;
      LAYER Metal3 ;
        RECT 424.27 12.00 424.93 12.66 ;
      LAYER Metal4 ;
        RECT 424.27 12.00 424.93 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 437.51 12.00 438.17 12.66 ;
      LAYER Metal6 ;
        RECT 437.51 12.00 438.17 12.66 ;
      LAYER Metal3 ;
        RECT 437.51 12.00 438.17 12.66 ;
      LAYER Metal4 ;
        RECT 437.51 12.00 438.17 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 466.83 12.00 467.49 12.66 ;
      LAYER Metal6 ;
        RECT 466.83 12.00 467.49 12.66 ;
      LAYER Metal3 ;
        RECT 466.83 12.00 467.49 12.66 ;
      LAYER Metal4 ;
        RECT 466.83 12.00 467.49 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.23 12.00 51.89 12.66 ;
      LAYER Metal6 ;
        RECT 51.23 12.00 51.89 12.66 ;
      LAYER Metal3 ;
        RECT 51.23 12.00 51.89 12.66 ;
      LAYER Metal4 ;
        RECT 51.23 12.00 51.89 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 480.07 12.00 480.73 12.66 ;
      LAYER Metal6 ;
        RECT 480.07 12.00 480.73 12.66 ;
      LAYER Metal3 ;
        RECT 480.07 12.00 480.73 12.66 ;
      LAYER Metal4 ;
        RECT 480.07 12.00 480.73 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 509.39 12.00 510.05 12.66 ;
      LAYER Metal6 ;
        RECT 509.39 12.00 510.05 12.66 ;
      LAYER Metal3 ;
        RECT 509.39 12.00 510.05 12.66 ;
      LAYER Metal4 ;
        RECT 509.39 12.00 510.05 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 522.63 12.00 523.29 12.66 ;
      LAYER Metal6 ;
        RECT 522.63 12.00 523.29 12.66 ;
      LAYER Metal3 ;
        RECT 522.63 12.00 523.29 12.66 ;
      LAYER Metal4 ;
        RECT 522.63 12.00 523.29 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 551.95 12.00 552.61 12.66 ;
      LAYER Metal6 ;
        RECT 551.95 12.00 552.61 12.66 ;
      LAYER Metal3 ;
        RECT 551.95 12.00 552.61 12.66 ;
      LAYER Metal4 ;
        RECT 551.95 12.00 552.61 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 565.19 12.00 565.85 12.66 ;
      LAYER Metal6 ;
        RECT 565.19 12.00 565.85 12.66 ;
      LAYER Metal3 ;
        RECT 565.19 12.00 565.85 12.66 ;
      LAYER Metal4 ;
        RECT 565.19 12.00 565.85 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 594.51 12.00 595.17 12.66 ;
      LAYER Metal6 ;
        RECT 594.51 12.00 595.17 12.66 ;
      LAYER Metal3 ;
        RECT 594.51 12.00 595.17 12.66 ;
      LAYER Metal4 ;
        RECT 594.51 12.00 595.17 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 607.75 12.00 608.41 12.66 ;
      LAYER Metal6 ;
        RECT 607.75 12.00 608.41 12.66 ;
      LAYER Metal3 ;
        RECT 607.75 12.00 608.41 12.66 ;
      LAYER Metal4 ;
        RECT 607.75 12.00 608.41 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 637.07 12.00 637.73 12.66 ;
      LAYER Metal6 ;
        RECT 637.07 12.00 637.73 12.66 ;
      LAYER Metal3 ;
        RECT 637.07 12.00 637.73 12.66 ;
      LAYER Metal4 ;
        RECT 637.07 12.00 637.73 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 650.31 12.00 650.97 12.66 ;
      LAYER Metal6 ;
        RECT 650.31 12.00 650.97 12.66 ;
      LAYER Metal3 ;
        RECT 650.31 12.00 650.97 12.66 ;
      LAYER Metal4 ;
        RECT 650.31 12.00 650.97 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 679.63 12.00 680.29 12.66 ;
      LAYER Metal6 ;
        RECT 679.63 12.00 680.29 12.66 ;
      LAYER Metal3 ;
        RECT 679.63 12.00 680.29 12.66 ;
      LAYER Metal4 ;
        RECT 679.63 12.00 680.29 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.47 12.00 65.13 12.66 ;
      LAYER Metal6 ;
        RECT 64.47 12.00 65.13 12.66 ;
      LAYER Metal3 ;
        RECT 64.47 12.00 65.13 12.66 ;
      LAYER Metal4 ;
        RECT 64.47 12.00 65.13 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 692.87 12.00 693.53 12.66 ;
      LAYER Metal6 ;
        RECT 692.87 12.00 693.53 12.66 ;
      LAYER Metal3 ;
        RECT 692.87 12.00 693.53 12.66 ;
      LAYER Metal4 ;
        RECT 692.87 12.00 693.53 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 722.19 12.00 722.85 12.66 ;
      LAYER Metal6 ;
        RECT 722.19 12.00 722.85 12.66 ;
      LAYER Metal3 ;
        RECT 722.19 12.00 722.85 12.66 ;
      LAYER Metal4 ;
        RECT 722.19 12.00 722.85 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.79 12.00 94.45 12.66 ;
      LAYER Metal6 ;
        RECT 93.79 12.00 94.45 12.66 ;
      LAYER Metal3 ;
        RECT 93.79 12.00 94.45 12.66 ;
      LAYER Metal4 ;
        RECT 93.79 12.00 94.45 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.03 12.00 107.69 12.66 ;
      LAYER Metal6 ;
        RECT 107.03 12.00 107.69 12.66 ;
      LAYER Metal3 ;
        RECT 107.03 12.00 107.69 12.66 ;
      LAYER Metal4 ;
        RECT 107.03 12.00 107.69 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.35 12.00 137.01 12.66 ;
      LAYER Metal6 ;
        RECT 136.35 12.00 137.01 12.66 ;
      LAYER Metal3 ;
        RECT 136.35 12.00 137.01 12.66 ;
      LAYER Metal4 ;
        RECT 136.35 12.00 137.01 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.59 12.00 150.25 12.66 ;
      LAYER Metal6 ;
        RECT 149.59 12.00 150.25 12.66 ;
      LAYER Metal3 ;
        RECT 149.59 12.00 150.25 12.66 ;
      LAYER Metal4 ;
        RECT 149.59 12.00 150.25 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.91 12.00 179.57 12.66 ;
      LAYER Metal6 ;
        RECT 178.91 12.00 179.57 12.66 ;
      LAYER Metal3 ;
        RECT 178.91 12.00 179.57 12.66 ;
      LAYER Metal4 ;
        RECT 178.91 12.00 179.57 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 192.15 12.00 192.81 12.66 ;
      LAYER Metal6 ;
        RECT 192.15 12.00 192.81 12.66 ;
      LAYER Metal3 ;
        RECT 192.15 12.00 192.81 12.66 ;
      LAYER Metal4 ;
        RECT 192.15 12.00 192.81 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.47 12.00 222.13 12.66 ;
      LAYER Metal6 ;
        RECT 221.47 12.00 222.13 12.66 ;
      LAYER Metal3 ;
        RECT 221.47 12.00 222.13 12.66 ;
      LAYER Metal4 ;
        RECT 221.47 12.00 222.13 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.95 12.00 30.61 12.66 ;
      LAYER Metal6 ;
        RECT 29.95 12.00 30.61 12.66 ;
      LAYER Metal3 ;
        RECT 29.95 12.00 30.61 12.66 ;
      LAYER Metal4 ;
        RECT 29.95 12.00 30.61 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.75 12.00 243.41 12.66 ;
      LAYER Metal6 ;
        RECT 242.75 12.00 243.41 12.66 ;
      LAYER Metal3 ;
        RECT 242.75 12.00 243.41 12.66 ;
      LAYER Metal4 ;
        RECT 242.75 12.00 243.41 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 255.99 12.00 256.65 12.66 ;
      LAYER Metal6 ;
        RECT 255.99 12.00 256.65 12.66 ;
      LAYER Metal3 ;
        RECT 255.99 12.00 256.65 12.66 ;
      LAYER Metal4 ;
        RECT 255.99 12.00 256.65 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.31 12.00 285.97 12.66 ;
      LAYER Metal6 ;
        RECT 285.31 12.00 285.97 12.66 ;
      LAYER Metal3 ;
        RECT 285.31 12.00 285.97 12.66 ;
      LAYER Metal4 ;
        RECT 285.31 12.00 285.97 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 298.55 12.00 299.21 12.66 ;
      LAYER Metal6 ;
        RECT 298.55 12.00 299.21 12.66 ;
      LAYER Metal3 ;
        RECT 298.55 12.00 299.21 12.66 ;
      LAYER Metal4 ;
        RECT 298.55 12.00 299.21 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 327.87 12.00 328.53 12.66 ;
      LAYER Metal6 ;
        RECT 327.87 12.00 328.53 12.66 ;
      LAYER Metal3 ;
        RECT 327.87 12.00 328.53 12.66 ;
      LAYER Metal4 ;
        RECT 327.87 12.00 328.53 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 341.11 12.00 341.77 12.66 ;
      LAYER Metal6 ;
        RECT 341.11 12.00 341.77 12.66 ;
      LAYER Metal3 ;
        RECT 341.11 12.00 341.77 12.66 ;
      LAYER Metal4 ;
        RECT 341.11 12.00 341.77 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 402.99 12.00 403.65 12.66 ;
      LAYER Metal6 ;
        RECT 402.99 12.00 403.65 12.66 ;
      LAYER Metal3 ;
        RECT 402.99 12.00 403.65 12.66 ;
      LAYER Metal4 ;
        RECT 402.99 12.00 403.65 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 416.23 12.00 416.89 12.66 ;
      LAYER Metal6 ;
        RECT 416.23 12.00 416.89 12.66 ;
      LAYER Metal3 ;
        RECT 416.23 12.00 416.89 12.66 ;
      LAYER Metal4 ;
        RECT 416.23 12.00 416.89 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 445.55 12.00 446.21 12.66 ;
      LAYER Metal6 ;
        RECT 445.55 12.00 446.21 12.66 ;
      LAYER Metal3 ;
        RECT 445.55 12.00 446.21 12.66 ;
      LAYER Metal4 ;
        RECT 445.55 12.00 446.21 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 458.79 12.00 459.45 12.66 ;
      LAYER Metal6 ;
        RECT 458.79 12.00 459.45 12.66 ;
      LAYER Metal3 ;
        RECT 458.79 12.00 459.45 12.66 ;
      LAYER Metal4 ;
        RECT 458.79 12.00 459.45 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.19 12.00 43.85 12.66 ;
      LAYER Metal6 ;
        RECT 43.19 12.00 43.85 12.66 ;
      LAYER Metal3 ;
        RECT 43.19 12.00 43.85 12.66 ;
      LAYER Metal4 ;
        RECT 43.19 12.00 43.85 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 488.11 12.00 488.77 12.66 ;
      LAYER Metal6 ;
        RECT 488.11 12.00 488.77 12.66 ;
      LAYER Metal3 ;
        RECT 488.11 12.00 488.77 12.66 ;
      LAYER Metal4 ;
        RECT 488.11 12.00 488.77 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 501.35 12.00 502.01 12.66 ;
      LAYER Metal6 ;
        RECT 501.35 12.00 502.01 12.66 ;
      LAYER Metal3 ;
        RECT 501.35 12.00 502.01 12.66 ;
      LAYER Metal4 ;
        RECT 501.35 12.00 502.01 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 530.67 12.00 531.33 12.66 ;
      LAYER Metal6 ;
        RECT 530.67 12.00 531.33 12.66 ;
      LAYER Metal3 ;
        RECT 530.67 12.00 531.33 12.66 ;
      LAYER Metal4 ;
        RECT 530.67 12.00 531.33 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 543.91 12.00 544.57 12.66 ;
      LAYER Metal6 ;
        RECT 543.91 12.00 544.57 12.66 ;
      LAYER Metal3 ;
        RECT 543.91 12.00 544.57 12.66 ;
      LAYER Metal4 ;
        RECT 543.91 12.00 544.57 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 573.23 12.00 573.89 12.66 ;
      LAYER Metal6 ;
        RECT 573.23 12.00 573.89 12.66 ;
      LAYER Metal3 ;
        RECT 573.23 12.00 573.89 12.66 ;
      LAYER Metal4 ;
        RECT 573.23 12.00 573.89 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 586.47 12.00 587.13 12.66 ;
      LAYER Metal6 ;
        RECT 586.47 12.00 587.13 12.66 ;
      LAYER Metal3 ;
        RECT 586.47 12.00 587.13 12.66 ;
      LAYER Metal4 ;
        RECT 586.47 12.00 587.13 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 615.79 12.00 616.45 12.66 ;
      LAYER Metal6 ;
        RECT 615.79 12.00 616.45 12.66 ;
      LAYER Metal3 ;
        RECT 615.79 12.00 616.45 12.66 ;
      LAYER Metal4 ;
        RECT 615.79 12.00 616.45 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 629.03 12.00 629.69 12.66 ;
      LAYER Metal6 ;
        RECT 629.03 12.00 629.69 12.66 ;
      LAYER Metal3 ;
        RECT 629.03 12.00 629.69 12.66 ;
      LAYER Metal4 ;
        RECT 629.03 12.00 629.69 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 658.35 12.00 659.01 12.66 ;
      LAYER Metal6 ;
        RECT 658.35 12.00 659.01 12.66 ;
      LAYER Metal3 ;
        RECT 658.35 12.00 659.01 12.66 ;
      LAYER Metal4 ;
        RECT 658.35 12.00 659.01 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 671.59 12.00 672.25 12.66 ;
      LAYER Metal6 ;
        RECT 671.59 12.00 672.25 12.66 ;
      LAYER Metal3 ;
        RECT 671.59 12.00 672.25 12.66 ;
      LAYER Metal4 ;
        RECT 671.59 12.00 672.25 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.51 12.00 73.17 12.66 ;
      LAYER Metal6 ;
        RECT 72.51 12.00 73.17 12.66 ;
      LAYER Metal3 ;
        RECT 72.51 12.00 73.17 12.66 ;
      LAYER Metal4 ;
        RECT 72.51 12.00 73.17 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 700.91 12.00 701.57 12.66 ;
      LAYER Metal6 ;
        RECT 700.91 12.00 701.57 12.66 ;
      LAYER Metal3 ;
        RECT 700.91 12.00 701.57 12.66 ;
      LAYER Metal4 ;
        RECT 700.91 12.00 701.57 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 714.15 12.00 714.81 12.66 ;
      LAYER Metal6 ;
        RECT 714.15 12.00 714.81 12.66 ;
      LAYER Metal3 ;
        RECT 714.15 12.00 714.81 12.66 ;
      LAYER Metal4 ;
        RECT 714.15 12.00 714.81 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.75 12.00 86.41 12.66 ;
      LAYER Metal6 ;
        RECT 85.75 12.00 86.41 12.66 ;
      LAYER Metal3 ;
        RECT 85.75 12.00 86.41 12.66 ;
      LAYER Metal4 ;
        RECT 85.75 12.00 86.41 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.07 12.00 115.73 12.66 ;
      LAYER Metal6 ;
        RECT 115.07 12.00 115.73 12.66 ;
      LAYER Metal3 ;
        RECT 115.07 12.00 115.73 12.66 ;
      LAYER Metal4 ;
        RECT 115.07 12.00 115.73 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.31 12.00 128.97 12.66 ;
      LAYER Metal6 ;
        RECT 128.31 12.00 128.97 12.66 ;
      LAYER Metal3 ;
        RECT 128.31 12.00 128.97 12.66 ;
      LAYER Metal4 ;
        RECT 128.31 12.00 128.97 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.63 12.00 158.29 12.66 ;
      LAYER Metal6 ;
        RECT 157.63 12.00 158.29 12.66 ;
      LAYER Metal3 ;
        RECT 157.63 12.00 158.29 12.66 ;
      LAYER Metal4 ;
        RECT 157.63 12.00 158.29 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 170.87 12.00 171.53 12.66 ;
      LAYER Metal6 ;
        RECT 170.87 12.00 171.53 12.66 ;
      LAYER Metal3 ;
        RECT 170.87 12.00 171.53 12.66 ;
      LAYER Metal4 ;
        RECT 170.87 12.00 171.53 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 200.19 12.00 200.85 12.66 ;
      LAYER Metal6 ;
        RECT 200.19 12.00 200.85 12.66 ;
      LAYER Metal3 ;
        RECT 200.19 12.00 200.85 12.66 ;
      LAYER Metal4 ;
        RECT 200.19 12.00 200.85 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 213.43 12.00 214.09 12.66 ;
      LAYER Metal6 ;
        RECT 213.43 12.00 214.09 12.66 ;
      LAYER Metal3 ;
        RECT 213.43 12.00 214.09 12.66 ;
      LAYER Metal4 ;
        RECT 213.43 12.00 214.09 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 24.49 12.00 25.15 12.66 ;
      LAYER Metal6 ;
        RECT 24.49 12.00 25.15 12.66 ;
      LAYER Metal3 ;
        RECT 24.49 12.00 25.15 12.66 ;
      LAYER Metal4 ;
        RECT 24.49 12.00 25.15 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 237.29 12.00 237.95 12.66 ;
      LAYER Metal6 ;
        RECT 237.29 12.00 237.95 12.66 ;
      LAYER Metal3 ;
        RECT 237.29 12.00 237.95 12.66 ;
      LAYER Metal4 ;
        RECT 237.29 12.00 237.95 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 261.45 12.00 262.11 12.66 ;
      LAYER Metal6 ;
        RECT 261.45 12.00 262.11 12.66 ;
      LAYER Metal3 ;
        RECT 261.45 12.00 262.11 12.66 ;
      LAYER Metal4 ;
        RECT 261.45 12.00 262.11 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 279.85 12.00 280.51 12.66 ;
      LAYER Metal6 ;
        RECT 279.85 12.00 280.51 12.66 ;
      LAYER Metal3 ;
        RECT 279.85 12.00 280.51 12.66 ;
      LAYER Metal4 ;
        RECT 279.85 12.00 280.51 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 304.01 12.00 304.67 12.66 ;
      LAYER Metal6 ;
        RECT 304.01 12.00 304.67 12.66 ;
      LAYER Metal3 ;
        RECT 304.01 12.00 304.67 12.66 ;
      LAYER Metal4 ;
        RECT 304.01 12.00 304.67 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 322.41 12.00 323.07 12.66 ;
      LAYER Metal6 ;
        RECT 322.41 12.00 323.07 12.66 ;
      LAYER Metal3 ;
        RECT 322.41 12.00 323.07 12.66 ;
      LAYER Metal4 ;
        RECT 322.41 12.00 323.07 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 346.57 12.00 347.23 12.66 ;
      LAYER Metal6 ;
        RECT 346.57 12.00 347.23 12.66 ;
      LAYER Metal3 ;
        RECT 346.57 12.00 347.23 12.66 ;
      LAYER Metal4 ;
        RECT 346.57 12.00 347.23 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 397.53 12.00 398.19 12.66 ;
      LAYER Metal6 ;
        RECT 397.53 12.00 398.19 12.66 ;
      LAYER Metal3 ;
        RECT 397.53 12.00 398.19 12.66 ;
      LAYER Metal4 ;
        RECT 397.53 12.00 398.19 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 421.69 12.00 422.35 12.66 ;
      LAYER Metal6 ;
        RECT 421.69 12.00 422.35 12.66 ;
      LAYER Metal3 ;
        RECT 421.69 12.00 422.35 12.66 ;
      LAYER Metal4 ;
        RECT 421.69 12.00 422.35 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 440.09 12.00 440.75 12.66 ;
      LAYER Metal6 ;
        RECT 440.09 12.00 440.75 12.66 ;
      LAYER Metal3 ;
        RECT 440.09 12.00 440.75 12.66 ;
      LAYER Metal4 ;
        RECT 440.09 12.00 440.75 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 464.25 12.00 464.91 12.66 ;
      LAYER Metal6 ;
        RECT 464.25 12.00 464.91 12.66 ;
      LAYER Metal3 ;
        RECT 464.25 12.00 464.91 12.66 ;
      LAYER Metal4 ;
        RECT 464.25 12.00 464.91 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 48.65 12.00 49.31 12.66 ;
      LAYER Metal6 ;
        RECT 48.65 12.00 49.31 12.66 ;
      LAYER Metal3 ;
        RECT 48.65 12.00 49.31 12.66 ;
      LAYER Metal4 ;
        RECT 48.65 12.00 49.31 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 482.65 12.00 483.31 12.66 ;
      LAYER Metal6 ;
        RECT 482.65 12.00 483.31 12.66 ;
      LAYER Metal3 ;
        RECT 482.65 12.00 483.31 12.66 ;
      LAYER Metal4 ;
        RECT 482.65 12.00 483.31 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 506.81 12.00 507.47 12.66 ;
      LAYER Metal6 ;
        RECT 506.81 12.00 507.47 12.66 ;
      LAYER Metal3 ;
        RECT 506.81 12.00 507.47 12.66 ;
      LAYER Metal4 ;
        RECT 506.81 12.00 507.47 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 525.21 12.00 525.87 12.66 ;
      LAYER Metal6 ;
        RECT 525.21 12.00 525.87 12.66 ;
      LAYER Metal3 ;
        RECT 525.21 12.00 525.87 12.66 ;
      LAYER Metal4 ;
        RECT 525.21 12.00 525.87 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 549.37 12.00 550.03 12.66 ;
      LAYER Metal6 ;
        RECT 549.37 12.00 550.03 12.66 ;
      LAYER Metal3 ;
        RECT 549.37 12.00 550.03 12.66 ;
      LAYER Metal4 ;
        RECT 549.37 12.00 550.03 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 567.77 12.00 568.43 12.66 ;
      LAYER Metal6 ;
        RECT 567.77 12.00 568.43 12.66 ;
      LAYER Metal3 ;
        RECT 567.77 12.00 568.43 12.66 ;
      LAYER Metal4 ;
        RECT 567.77 12.00 568.43 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 591.93 12.00 592.59 12.66 ;
      LAYER Metal6 ;
        RECT 591.93 12.00 592.59 12.66 ;
      LAYER Metal3 ;
        RECT 591.93 12.00 592.59 12.66 ;
      LAYER Metal4 ;
        RECT 591.93 12.00 592.59 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 610.33 12.00 610.99 12.66 ;
      LAYER Metal6 ;
        RECT 610.33 12.00 610.99 12.66 ;
      LAYER Metal3 ;
        RECT 610.33 12.00 610.99 12.66 ;
      LAYER Metal4 ;
        RECT 610.33 12.00 610.99 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 634.49 12.00 635.15 12.66 ;
      LAYER Metal6 ;
        RECT 634.49 12.00 635.15 12.66 ;
      LAYER Metal3 ;
        RECT 634.49 12.00 635.15 12.66 ;
      LAYER Metal4 ;
        RECT 634.49 12.00 635.15 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 652.89 12.00 653.55 12.66 ;
      LAYER Metal6 ;
        RECT 652.89 12.00 653.55 12.66 ;
      LAYER Metal3 ;
        RECT 652.89 12.00 653.55 12.66 ;
      LAYER Metal4 ;
        RECT 652.89 12.00 653.55 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 677.05 12.00 677.71 12.66 ;
      LAYER Metal6 ;
        RECT 677.05 12.00 677.71 12.66 ;
      LAYER Metal3 ;
        RECT 677.05 12.00 677.71 12.66 ;
      LAYER Metal4 ;
        RECT 677.05 12.00 677.71 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.05 12.00 67.71 12.66 ;
      LAYER Metal6 ;
        RECT 67.05 12.00 67.71 12.66 ;
      LAYER Metal3 ;
        RECT 67.05 12.00 67.71 12.66 ;
      LAYER Metal4 ;
        RECT 67.05 12.00 67.71 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 695.45 12.00 696.11 12.66 ;
      LAYER Metal6 ;
        RECT 695.45 12.00 696.11 12.66 ;
      LAYER Metal3 ;
        RECT 695.45 12.00 696.11 12.66 ;
      LAYER Metal4 ;
        RECT 695.45 12.00 696.11 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 719.61 12.00 720.27 12.66 ;
      LAYER Metal6 ;
        RECT 719.61 12.00 720.27 12.66 ;
      LAYER Metal3 ;
        RECT 719.61 12.00 720.27 12.66 ;
      LAYER Metal4 ;
        RECT 719.61 12.00 720.27 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 91.21 12.00 91.87 12.66 ;
      LAYER Metal6 ;
        RECT 91.21 12.00 91.87 12.66 ;
      LAYER Metal3 ;
        RECT 91.21 12.00 91.87 12.66 ;
      LAYER Metal4 ;
        RECT 91.21 12.00 91.87 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 109.61 12.00 110.27 12.66 ;
      LAYER Metal6 ;
        RECT 109.61 12.00 110.27 12.66 ;
      LAYER Metal3 ;
        RECT 109.61 12.00 110.27 12.66 ;
      LAYER Metal4 ;
        RECT 109.61 12.00 110.27 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 133.77 12.00 134.43 12.66 ;
      LAYER Metal6 ;
        RECT 133.77 12.00 134.43 12.66 ;
      LAYER Metal3 ;
        RECT 133.77 12.00 134.43 12.66 ;
      LAYER Metal4 ;
        RECT 133.77 12.00 134.43 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 152.17 12.00 152.83 12.66 ;
      LAYER Metal6 ;
        RECT 152.17 12.00 152.83 12.66 ;
      LAYER Metal3 ;
        RECT 152.17 12.00 152.83 12.66 ;
      LAYER Metal4 ;
        RECT 152.17 12.00 152.83 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 176.33 12.00 176.99 12.66 ;
      LAYER Metal6 ;
        RECT 176.33 12.00 176.99 12.66 ;
      LAYER Metal3 ;
        RECT 176.33 12.00 176.99 12.66 ;
      LAYER Metal4 ;
        RECT 176.33 12.00 176.99 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 194.73 12.00 195.39 12.66 ;
      LAYER Metal6 ;
        RECT 194.73 12.00 195.39 12.66 ;
      LAYER Metal3 ;
        RECT 194.73 12.00 195.39 12.66 ;
      LAYER Metal4 ;
        RECT 194.73 12.00 195.39 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.89 12.00 219.55 12.66 ;
      LAYER Metal6 ;
        RECT 218.89 12.00 219.55 12.66 ;
      LAYER Metal3 ;
        RECT 218.89 12.00 219.55 12.66 ;
      LAYER Metal4 ;
        RECT 218.89 12.00 219.55 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 27.37 12.00 28.03 12.66 ;
      LAYER Metal6 ;
        RECT 27.37 12.00 28.03 12.66 ;
      LAYER Metal3 ;
        RECT 27.37 12.00 28.03 12.66 ;
      LAYER Metal4 ;
        RECT 27.37 12.00 28.03 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 240.17 12.00 240.83 12.66 ;
      LAYER Metal6 ;
        RECT 240.17 12.00 240.83 12.66 ;
      LAYER Metal3 ;
        RECT 240.17 12.00 240.83 12.66 ;
      LAYER Metal4 ;
        RECT 240.17 12.00 240.83 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 258.57 12.00 259.23 12.66 ;
      LAYER Metal6 ;
        RECT 258.57 12.00 259.23 12.66 ;
      LAYER Metal3 ;
        RECT 258.57 12.00 259.23 12.66 ;
      LAYER Metal4 ;
        RECT 258.57 12.00 259.23 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 282.73 12.00 283.39 12.66 ;
      LAYER Metal6 ;
        RECT 282.73 12.00 283.39 12.66 ;
      LAYER Metal3 ;
        RECT 282.73 12.00 283.39 12.66 ;
      LAYER Metal4 ;
        RECT 282.73 12.00 283.39 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 301.13 12.00 301.79 12.66 ;
      LAYER Metal6 ;
        RECT 301.13 12.00 301.79 12.66 ;
      LAYER Metal3 ;
        RECT 301.13 12.00 301.79 12.66 ;
      LAYER Metal4 ;
        RECT 301.13 12.00 301.79 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 325.29 12.00 325.95 12.66 ;
      LAYER Metal6 ;
        RECT 325.29 12.00 325.95 12.66 ;
      LAYER Metal3 ;
        RECT 325.29 12.00 325.95 12.66 ;
      LAYER Metal4 ;
        RECT 325.29 12.00 325.95 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 343.69 12.00 344.35 12.66 ;
      LAYER Metal6 ;
        RECT 343.69 12.00 344.35 12.66 ;
      LAYER Metal3 ;
        RECT 343.69 12.00 344.35 12.66 ;
      LAYER Metal4 ;
        RECT 343.69 12.00 344.35 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 400.41 12.00 401.07 12.66 ;
      LAYER Metal6 ;
        RECT 400.41 12.00 401.07 12.66 ;
      LAYER Metal3 ;
        RECT 400.41 12.00 401.07 12.66 ;
      LAYER Metal4 ;
        RECT 400.41 12.00 401.07 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 418.81 12.00 419.47 12.66 ;
      LAYER Metal6 ;
        RECT 418.81 12.00 419.47 12.66 ;
      LAYER Metal3 ;
        RECT 418.81 12.00 419.47 12.66 ;
      LAYER Metal4 ;
        RECT 418.81 12.00 419.47 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 442.97 12.00 443.63 12.66 ;
      LAYER Metal6 ;
        RECT 442.97 12.00 443.63 12.66 ;
      LAYER Metal3 ;
        RECT 442.97 12.00 443.63 12.66 ;
      LAYER Metal4 ;
        RECT 442.97 12.00 443.63 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 461.37 12.00 462.03 12.66 ;
      LAYER Metal6 ;
        RECT 461.37 12.00 462.03 12.66 ;
      LAYER Metal3 ;
        RECT 461.37 12.00 462.03 12.66 ;
      LAYER Metal4 ;
        RECT 461.37 12.00 462.03 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 45.77 12.00 46.43 12.66 ;
      LAYER Metal6 ;
        RECT 45.77 12.00 46.43 12.66 ;
      LAYER Metal3 ;
        RECT 45.77 12.00 46.43 12.66 ;
      LAYER Metal4 ;
        RECT 45.77 12.00 46.43 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 485.53 12.00 486.19 12.66 ;
      LAYER Metal6 ;
        RECT 485.53 12.00 486.19 12.66 ;
      LAYER Metal3 ;
        RECT 485.53 12.00 486.19 12.66 ;
      LAYER Metal4 ;
        RECT 485.53 12.00 486.19 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 503.93 12.00 504.59 12.66 ;
      LAYER Metal6 ;
        RECT 503.93 12.00 504.59 12.66 ;
      LAYER Metal3 ;
        RECT 503.93 12.00 504.59 12.66 ;
      LAYER Metal4 ;
        RECT 503.93 12.00 504.59 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 528.09 12.00 528.75 12.66 ;
      LAYER Metal6 ;
        RECT 528.09 12.00 528.75 12.66 ;
      LAYER Metal3 ;
        RECT 528.09 12.00 528.75 12.66 ;
      LAYER Metal4 ;
        RECT 528.09 12.00 528.75 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 546.49 12.00 547.15 12.66 ;
      LAYER Metal6 ;
        RECT 546.49 12.00 547.15 12.66 ;
      LAYER Metal3 ;
        RECT 546.49 12.00 547.15 12.66 ;
      LAYER Metal4 ;
        RECT 546.49 12.00 547.15 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 570.65 12.00 571.31 12.66 ;
      LAYER Metal6 ;
        RECT 570.65 12.00 571.31 12.66 ;
      LAYER Metal3 ;
        RECT 570.65 12.00 571.31 12.66 ;
      LAYER Metal4 ;
        RECT 570.65 12.00 571.31 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 589.05 12.00 589.71 12.66 ;
      LAYER Metal6 ;
        RECT 589.05 12.00 589.71 12.66 ;
      LAYER Metal3 ;
        RECT 589.05 12.00 589.71 12.66 ;
      LAYER Metal4 ;
        RECT 589.05 12.00 589.71 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 613.21 12.00 613.87 12.66 ;
      LAYER Metal6 ;
        RECT 613.21 12.00 613.87 12.66 ;
      LAYER Metal3 ;
        RECT 613.21 12.00 613.87 12.66 ;
      LAYER Metal4 ;
        RECT 613.21 12.00 613.87 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 631.61 12.00 632.27 12.66 ;
      LAYER Metal6 ;
        RECT 631.61 12.00 632.27 12.66 ;
      LAYER Metal3 ;
        RECT 631.61 12.00 632.27 12.66 ;
      LAYER Metal4 ;
        RECT 631.61 12.00 632.27 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 655.77 12.00 656.43 12.66 ;
      LAYER Metal6 ;
        RECT 655.77 12.00 656.43 12.66 ;
      LAYER Metal3 ;
        RECT 655.77 12.00 656.43 12.66 ;
      LAYER Metal4 ;
        RECT 655.77 12.00 656.43 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 674.17 12.00 674.83 12.66 ;
      LAYER Metal6 ;
        RECT 674.17 12.00 674.83 12.66 ;
      LAYER Metal3 ;
        RECT 674.17 12.00 674.83 12.66 ;
      LAYER Metal4 ;
        RECT 674.17 12.00 674.83 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.93 12.00 70.59 12.66 ;
      LAYER Metal6 ;
        RECT 69.93 12.00 70.59 12.66 ;
      LAYER Metal3 ;
        RECT 69.93 12.00 70.59 12.66 ;
      LAYER Metal4 ;
        RECT 69.93 12.00 70.59 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 698.33 12.00 698.99 12.66 ;
      LAYER Metal6 ;
        RECT 698.33 12.00 698.99 12.66 ;
      LAYER Metal3 ;
        RECT 698.33 12.00 698.99 12.66 ;
      LAYER Metal4 ;
        RECT 698.33 12.00 698.99 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 716.73 12.00 717.39 12.66 ;
      LAYER Metal6 ;
        RECT 716.73 12.00 717.39 12.66 ;
      LAYER Metal3 ;
        RECT 716.73 12.00 717.39 12.66 ;
      LAYER Metal4 ;
        RECT 716.73 12.00 717.39 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 88.33 12.00 88.99 12.66 ;
      LAYER Metal6 ;
        RECT 88.33 12.00 88.99 12.66 ;
      LAYER Metal3 ;
        RECT 88.33 12.00 88.99 12.66 ;
      LAYER Metal4 ;
        RECT 88.33 12.00 88.99 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 112.49 12.00 113.15 12.66 ;
      LAYER Metal6 ;
        RECT 112.49 12.00 113.15 12.66 ;
      LAYER Metal3 ;
        RECT 112.49 12.00 113.15 12.66 ;
      LAYER Metal4 ;
        RECT 112.49 12.00 113.15 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 130.89 12.00 131.55 12.66 ;
      LAYER Metal6 ;
        RECT 130.89 12.00 131.55 12.66 ;
      LAYER Metal3 ;
        RECT 130.89 12.00 131.55 12.66 ;
      LAYER Metal4 ;
        RECT 130.89 12.00 131.55 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 155.05 12.00 155.71 12.66 ;
      LAYER Metal6 ;
        RECT 155.05 12.00 155.71 12.66 ;
      LAYER Metal3 ;
        RECT 155.05 12.00 155.71 12.66 ;
      LAYER Metal4 ;
        RECT 155.05 12.00 155.71 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 173.45 12.00 174.11 12.66 ;
      LAYER Metal6 ;
        RECT 173.45 12.00 174.11 12.66 ;
      LAYER Metal3 ;
        RECT 173.45 12.00 174.11 12.66 ;
      LAYER Metal4 ;
        RECT 173.45 12.00 174.11 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 197.61 12.00 198.27 12.66 ;
      LAYER Metal6 ;
        RECT 197.61 12.00 198.27 12.66 ;
      LAYER Metal3 ;
        RECT 197.61 12.00 198.27 12.66 ;
      LAYER Metal4 ;
        RECT 197.61 12.00 198.27 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 216.01 12.00 216.67 12.66 ;
      LAYER Metal6 ;
        RECT 216.01 12.00 216.67 12.66 ;
      LAYER Metal3 ;
        RECT 216.01 12.00 216.67 12.66 ;
      LAYER Metal4 ;
        RECT 216.01 12.00 216.67 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 379.9 12.00 380.56 12.66 ;
      LAYER Metal6 ;
        RECT 379.9 12.00 380.56 12.66 ;
      LAYER Metal3 ;
        RECT 379.9 12.00 380.56 12.66 ;
      LAYER Metal4 ;
        RECT 379.9 12.00 380.56 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 364.2 12.00 364.86 12.66 ;
      LAYER Metal6 ;
        RECT 364.2 12.00 364.86 12.66 ;
      LAYER Metal3 ;
        RECT 364.2 12.00 364.86 12.66 ;
      LAYER Metal4 ;
        RECT 364.2 12.00 364.86 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 202.2 763.02 207.2 ;
        RECT 0 0 763.02 5 ;
      LAYER Metal2 ;
        RECT 758.02 0 763.02 207.2 ;
        RECT 0 0 5 207.2 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 196.6 757.42 201.6 ;
        RECT 5.6 5.6 757.42 10.6 ;
      LAYER Metal2 ;
        RECT 752.42 5.6 757.42 201.6 ;
        RECT 5.6 5.6 10.6 201.6 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 751.015 195.24 ;
    LAYER Metal2 ;
      RECT 12 12 751.015 195.24 ;
    LAYER Metal3 ;
      RECT 12 12 751.015 195.24 ;
    LAYER Metal4 ;
      RECT 12 12 751.015 195.24 ;
    LAYER Metal5 ;
      RECT 12 12 751.015 195.24 ;
    LAYER Metal6 ;
      RECT 12 12 751.015 195.24 ;
  END
END MEM2_512X32

END LIBRARY
