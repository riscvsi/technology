VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MEM2_2048X32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2_2048X32 0 0 ;
  SIZE 761.745 BY 522.75 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 303.625 12.66 304.285 ;
      LAYER Metal6 ;
        RECT 12 303.625 12.66 304.285 ;
      LAYER Metal3 ;
        RECT 12 303.625 12.66 304.285 ;
      LAYER Metal4 ;
        RECT 12 303.625 12.66 304.285 ;
    END
  END A1[0]
  PIN A1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 260.785 12.66 261.445 ;
      LAYER Metal6 ;
        RECT 12 260.785 12.66 261.445 ;
      LAYER Metal3 ;
        RECT 12 260.785 12.66 261.445 ;
      LAYER Metal4 ;
        RECT 12 260.785 12.66 261.445 ;
    END
  END A1[10]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 297.505 12.66 298.165 ;
      LAYER Metal6 ;
        RECT 12 297.505 12.66 298.165 ;
      LAYER Metal3 ;
        RECT 12 297.505 12.66 298.165 ;
      LAYER Metal4 ;
        RECT 12 297.505 12.66 298.165 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 294.405 12.66 295.065 ;
      LAYER Metal6 ;
        RECT 12 294.405 12.66 295.065 ;
      LAYER Metal3 ;
        RECT 12 294.405 12.66 295.065 ;
      LAYER Metal4 ;
        RECT 12 294.405 12.66 295.065 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 288.285 12.66 288.945 ;
      LAYER Metal6 ;
        RECT 12 288.285 12.66 288.945 ;
      LAYER Metal3 ;
        RECT 12 288.285 12.66 288.945 ;
      LAYER Metal4 ;
        RECT 12 288.285 12.66 288.945 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 285.265 12.66 285.925 ;
      LAYER Metal6 ;
        RECT 12 285.265 12.66 285.925 ;
      LAYER Metal3 ;
        RECT 12 285.265 12.66 285.925 ;
      LAYER Metal4 ;
        RECT 12 285.265 12.66 285.925 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 282.165 12.66 282.825 ;
      LAYER Metal6 ;
        RECT 12 282.165 12.66 282.825 ;
      LAYER Metal3 ;
        RECT 12 282.165 12.66 282.825 ;
      LAYER Metal4 ;
        RECT 12 282.165 12.66 282.825 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 276.045 12.66 276.705 ;
      LAYER Metal6 ;
        RECT 12 276.045 12.66 276.705 ;
      LAYER Metal3 ;
        RECT 12 276.045 12.66 276.705 ;
      LAYER Metal4 ;
        RECT 12 276.045 12.66 276.705 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 273.025 12.66 273.685 ;
      LAYER Metal6 ;
        RECT 12 273.025 12.66 273.685 ;
      LAYER Metal3 ;
        RECT 12 273.025 12.66 273.685 ;
      LAYER Metal4 ;
        RECT 12 273.025 12.66 273.685 ;
    END
  END A1[7]
  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 269.925 12.66 270.585 ;
      LAYER Metal6 ;
        RECT 12 269.925 12.66 270.585 ;
      LAYER Metal3 ;
        RECT 12 269.925 12.66 270.585 ;
      LAYER Metal4 ;
        RECT 12 269.925 12.66 270.585 ;
    END
  END A1[8]
  PIN A1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 263.805 12.66 264.465 ;
      LAYER Metal6 ;
        RECT 12 263.805 12.66 264.465 ;
      LAYER Metal3 ;
        RECT 12 263.805 12.66 264.465 ;
      LAYER Metal4 ;
        RECT 12 263.805 12.66 264.465 ;
    END
  END A1[9]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 213.125 12.66 213.785 ;
      LAYER Metal6 ;
        RECT 12 213.125 12.66 213.785 ;
      LAYER Metal3 ;
        RECT 12 213.125 12.66 213.785 ;
      LAYER Metal4 ;
        RECT 12 213.125 12.66 213.785 ;
    END
  END A2[0]
  PIN A2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 255.965 12.66 256.625 ;
      LAYER Metal6 ;
        RECT 12 255.965 12.66 256.625 ;
      LAYER Metal3 ;
        RECT 12 255.965 12.66 256.625 ;
      LAYER Metal4 ;
        RECT 12 255.965 12.66 256.625 ;
    END
  END A2[10]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 219.245 12.66 219.905 ;
      LAYER Metal6 ;
        RECT 12 219.245 12.66 219.905 ;
      LAYER Metal3 ;
        RECT 12 219.245 12.66 219.905 ;
      LAYER Metal4 ;
        RECT 12 219.245 12.66 219.905 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 222.345 12.66 223.005 ;
      LAYER Metal6 ;
        RECT 12 222.345 12.66 223.005 ;
      LAYER Metal3 ;
        RECT 12 222.345 12.66 223.005 ;
      LAYER Metal4 ;
        RECT 12 222.345 12.66 223.005 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 228.465 12.66 229.125 ;
      LAYER Metal6 ;
        RECT 12 228.465 12.66 229.125 ;
      LAYER Metal3 ;
        RECT 12 228.465 12.66 229.125 ;
      LAYER Metal4 ;
        RECT 12 228.465 12.66 229.125 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 231.485 12.66 232.145 ;
      LAYER Metal6 ;
        RECT 12 231.485 12.66 232.145 ;
      LAYER Metal3 ;
        RECT 12 231.485 12.66 232.145 ;
      LAYER Metal4 ;
        RECT 12 231.485 12.66 232.145 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 234.585 12.66 235.245 ;
      LAYER Metal6 ;
        RECT 12 234.585 12.66 235.245 ;
      LAYER Metal3 ;
        RECT 12 234.585 12.66 235.245 ;
      LAYER Metal4 ;
        RECT 12 234.585 12.66 235.245 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 240.705 12.66 241.365 ;
      LAYER Metal6 ;
        RECT 12 240.705 12.66 241.365 ;
      LAYER Metal3 ;
        RECT 12 240.705 12.66 241.365 ;
      LAYER Metal4 ;
        RECT 12 240.705 12.66 241.365 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 243.725 12.66 244.385 ;
      LAYER Metal6 ;
        RECT 12 243.725 12.66 244.385 ;
      LAYER Metal3 ;
        RECT 12 243.725 12.66 244.385 ;
      LAYER Metal4 ;
        RECT 12 243.725 12.66 244.385 ;
    END
  END A2[7]
  PIN A2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 246.825 12.66 247.485 ;
      LAYER Metal6 ;
        RECT 12 246.825 12.66 247.485 ;
      LAYER Metal3 ;
        RECT 12 246.825 12.66 247.485 ;
      LAYER Metal4 ;
        RECT 12 246.825 12.66 247.485 ;
    END
  END A2[8]
  PIN A2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 252.945 12.66 253.605 ;
      LAYER Metal6 ;
        RECT 12 252.945 12.66 253.605 ;
      LAYER Metal3 ;
        RECT 12 252.945 12.66 253.605 ;
      LAYER Metal4 ;
        RECT 12 252.945 12.66 253.605 ;
    END
  END A2[9]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 373.61 12 374.27 12.66 ;
      LAYER Metal6 ;
        RECT 373.61 12 374.27 12.66 ;
      LAYER Metal3 ;
        RECT 373.61 12 374.27 12.66 ;
      LAYER Metal4 ;
        RECT 373.61 12 374.27 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.6 12 367.26 12.66 ;
      LAYER Metal6 ;
        RECT 366.6 12 367.26 12.66 ;
      LAYER Metal3 ;
        RECT 366.6 12 367.26 12.66 ;
      LAYER Metal4 ;
        RECT 366.6 12 367.26 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 382.235 12 382.895 12.66 ;
      LAYER Metal6 ;
        RECT 382.235 12 382.895 12.66 ;
      LAYER Metal3 ;
        RECT 382.235 12 382.895 12.66 ;
      LAYER Metal4 ;
        RECT 382.235 12 382.895 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 357.975 12 358.635 12.66 ;
      LAYER Metal6 ;
        RECT 357.975 12 358.635 12.66 ;
      LAYER Metal3 ;
        RECT 357.975 12 358.635 12.66 ;
      LAYER Metal4 ;
        RECT 357.975 12 358.635 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 21.91 12 22.57 12.66 ;
      LAYER Metal6 ;
        RECT 21.91 12 22.57 12.66 ;
      LAYER Metal3 ;
        RECT 21.91 12 22.57 12.66 ;
      LAYER Metal4 ;
        RECT 21.91 12 22.57 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.71 12 235.37 12.66 ;
      LAYER Metal6 ;
        RECT 234.71 12 235.37 12.66 ;
      LAYER Metal3 ;
        RECT 234.71 12 235.37 12.66 ;
      LAYER Metal4 ;
        RECT 234.71 12 235.37 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.03 12 264.69 12.66 ;
      LAYER Metal6 ;
        RECT 264.03 12 264.69 12.66 ;
      LAYER Metal3 ;
        RECT 264.03 12 264.69 12.66 ;
      LAYER Metal4 ;
        RECT 264.03 12 264.69 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 277.27 12 277.93 12.66 ;
      LAYER Metal6 ;
        RECT 277.27 12 277.93 12.66 ;
      LAYER Metal3 ;
        RECT 277.27 12 277.93 12.66 ;
      LAYER Metal4 ;
        RECT 277.27 12 277.93 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.59 12 307.25 12.66 ;
      LAYER Metal6 ;
        RECT 306.59 12 307.25 12.66 ;
      LAYER Metal3 ;
        RECT 306.59 12 307.25 12.66 ;
      LAYER Metal4 ;
        RECT 306.59 12 307.25 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 319.83 12 320.49 12.66 ;
      LAYER Metal6 ;
        RECT 319.83 12 320.49 12.66 ;
      LAYER Metal3 ;
        RECT 319.83 12 320.49 12.66 ;
      LAYER Metal4 ;
        RECT 319.83 12 320.49 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.15 12 349.81 12.66 ;
      LAYER Metal6 ;
        RECT 349.15 12 349.81 12.66 ;
      LAYER Metal3 ;
        RECT 349.15 12 349.81 12.66 ;
      LAYER Metal4 ;
        RECT 349.15 12 349.81 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 391.06 12 391.72 12.66 ;
      LAYER Metal6 ;
        RECT 391.06 12 391.72 12.66 ;
      LAYER Metal3 ;
        RECT 391.06 12 391.72 12.66 ;
      LAYER Metal4 ;
        RECT 391.06 12 391.72 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 420.38 12 421.04 12.66 ;
      LAYER Metal6 ;
        RECT 420.38 12 421.04 12.66 ;
      LAYER Metal3 ;
        RECT 420.38 12 421.04 12.66 ;
      LAYER Metal4 ;
        RECT 420.38 12 421.04 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 433.62 12 434.28 12.66 ;
      LAYER Metal6 ;
        RECT 433.62 12 434.28 12.66 ;
      LAYER Metal3 ;
        RECT 433.62 12 434.28 12.66 ;
      LAYER Metal4 ;
        RECT 433.62 12 434.28 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 462.94 12 463.6 12.66 ;
      LAYER Metal6 ;
        RECT 462.94 12 463.6 12.66 ;
      LAYER Metal3 ;
        RECT 462.94 12 463.6 12.66 ;
      LAYER Metal4 ;
        RECT 462.94 12 463.6 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.23 12 51.89 12.66 ;
      LAYER Metal6 ;
        RECT 51.23 12 51.89 12.66 ;
      LAYER Metal3 ;
        RECT 51.23 12 51.89 12.66 ;
      LAYER Metal4 ;
        RECT 51.23 12 51.89 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 476.18 12 476.84 12.66 ;
      LAYER Metal6 ;
        RECT 476.18 12 476.84 12.66 ;
      LAYER Metal3 ;
        RECT 476.18 12 476.84 12.66 ;
      LAYER Metal4 ;
        RECT 476.18 12 476.84 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 505.5 12 506.16 12.66 ;
      LAYER Metal6 ;
        RECT 505.5 12 506.16 12.66 ;
      LAYER Metal3 ;
        RECT 505.5 12 506.16 12.66 ;
      LAYER Metal4 ;
        RECT 505.5 12 506.16 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 518.74 12 519.4 12.66 ;
      LAYER Metal6 ;
        RECT 518.74 12 519.4 12.66 ;
      LAYER Metal3 ;
        RECT 518.74 12 519.4 12.66 ;
      LAYER Metal4 ;
        RECT 518.74 12 519.4 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 548.06 12 548.72 12.66 ;
      LAYER Metal6 ;
        RECT 548.06 12 548.72 12.66 ;
      LAYER Metal3 ;
        RECT 548.06 12 548.72 12.66 ;
      LAYER Metal4 ;
        RECT 548.06 12 548.72 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 561.3 12 561.96 12.66 ;
      LAYER Metal6 ;
        RECT 561.3 12 561.96 12.66 ;
      LAYER Metal3 ;
        RECT 561.3 12 561.96 12.66 ;
      LAYER Metal4 ;
        RECT 561.3 12 561.96 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 590.62 12 591.28 12.66 ;
      LAYER Metal6 ;
        RECT 590.62 12 591.28 12.66 ;
      LAYER Metal3 ;
        RECT 590.62 12 591.28 12.66 ;
      LAYER Metal4 ;
        RECT 590.62 12 591.28 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 603.86 12 604.52 12.66 ;
      LAYER Metal6 ;
        RECT 603.86 12 604.52 12.66 ;
      LAYER Metal3 ;
        RECT 603.86 12 604.52 12.66 ;
      LAYER Metal4 ;
        RECT 603.86 12 604.52 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 633.18 12 633.84 12.66 ;
      LAYER Metal6 ;
        RECT 633.18 12 633.84 12.66 ;
      LAYER Metal3 ;
        RECT 633.18 12 633.84 12.66 ;
      LAYER Metal4 ;
        RECT 633.18 12 633.84 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 646.42 12 647.08 12.66 ;
      LAYER Metal6 ;
        RECT 646.42 12 647.08 12.66 ;
      LAYER Metal3 ;
        RECT 646.42 12 647.08 12.66 ;
      LAYER Metal4 ;
        RECT 646.42 12 647.08 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 675.74 12 676.4 12.66 ;
      LAYER Metal6 ;
        RECT 675.74 12 676.4 12.66 ;
      LAYER Metal3 ;
        RECT 675.74 12 676.4 12.66 ;
      LAYER Metal4 ;
        RECT 675.74 12 676.4 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.47 12 65.13 12.66 ;
      LAYER Metal6 ;
        RECT 64.47 12 65.13 12.66 ;
      LAYER Metal3 ;
        RECT 64.47 12 65.13 12.66 ;
      LAYER Metal4 ;
        RECT 64.47 12 65.13 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 688.98 12 689.64 12.66 ;
      LAYER Metal6 ;
        RECT 688.98 12 689.64 12.66 ;
      LAYER Metal3 ;
        RECT 688.98 12 689.64 12.66 ;
      LAYER Metal4 ;
        RECT 688.98 12 689.64 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 718.3 12 718.96 12.66 ;
      LAYER Metal6 ;
        RECT 718.3 12 718.96 12.66 ;
      LAYER Metal3 ;
        RECT 718.3 12 718.96 12.66 ;
      LAYER Metal4 ;
        RECT 718.3 12 718.96 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.79 12 94.45 12.66 ;
      LAYER Metal6 ;
        RECT 93.79 12 94.45 12.66 ;
      LAYER Metal3 ;
        RECT 93.79 12 94.45 12.66 ;
      LAYER Metal4 ;
        RECT 93.79 12 94.45 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.03 12 107.69 12.66 ;
      LAYER Metal6 ;
        RECT 107.03 12 107.69 12.66 ;
      LAYER Metal3 ;
        RECT 107.03 12 107.69 12.66 ;
      LAYER Metal4 ;
        RECT 107.03 12 107.69 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.35 12 137.01 12.66 ;
      LAYER Metal6 ;
        RECT 136.35 12 137.01 12.66 ;
      LAYER Metal3 ;
        RECT 136.35 12 137.01 12.66 ;
      LAYER Metal4 ;
        RECT 136.35 12 137.01 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.59 12 150.25 12.66 ;
      LAYER Metal6 ;
        RECT 149.59 12 150.25 12.66 ;
      LAYER Metal3 ;
        RECT 149.59 12 150.25 12.66 ;
      LAYER Metal4 ;
        RECT 149.59 12 150.25 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.91 12 179.57 12.66 ;
      LAYER Metal6 ;
        RECT 178.91 12 179.57 12.66 ;
      LAYER Metal3 ;
        RECT 178.91 12 179.57 12.66 ;
      LAYER Metal4 ;
        RECT 178.91 12 179.57 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 192.15 12 192.81 12.66 ;
      LAYER Metal6 ;
        RECT 192.15 12 192.81 12.66 ;
      LAYER Metal3 ;
        RECT 192.15 12 192.81 12.66 ;
      LAYER Metal4 ;
        RECT 192.15 12 192.81 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.47 12 222.13 12.66 ;
      LAYER Metal6 ;
        RECT 221.47 12 222.13 12.66 ;
      LAYER Metal3 ;
        RECT 221.47 12 222.13 12.66 ;
      LAYER Metal4 ;
        RECT 221.47 12 222.13 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.95 12 30.61 12.66 ;
      LAYER Metal6 ;
        RECT 29.95 12 30.61 12.66 ;
      LAYER Metal3 ;
        RECT 29.95 12 30.61 12.66 ;
      LAYER Metal4 ;
        RECT 29.95 12 30.61 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.75 12 243.41 12.66 ;
      LAYER Metal6 ;
        RECT 242.75 12 243.41 12.66 ;
      LAYER Metal3 ;
        RECT 242.75 12 243.41 12.66 ;
      LAYER Metal4 ;
        RECT 242.75 12 243.41 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 255.99 12 256.65 12.66 ;
      LAYER Metal6 ;
        RECT 255.99 12 256.65 12.66 ;
      LAYER Metal3 ;
        RECT 255.99 12 256.65 12.66 ;
      LAYER Metal4 ;
        RECT 255.99 12 256.65 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.31 12 285.97 12.66 ;
      LAYER Metal6 ;
        RECT 285.31 12 285.97 12.66 ;
      LAYER Metal3 ;
        RECT 285.31 12 285.97 12.66 ;
      LAYER Metal4 ;
        RECT 285.31 12 285.97 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 298.55 12 299.21 12.66 ;
      LAYER Metal6 ;
        RECT 298.55 12 299.21 12.66 ;
      LAYER Metal3 ;
        RECT 298.55 12 299.21 12.66 ;
      LAYER Metal4 ;
        RECT 298.55 12 299.21 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 327.87 12 328.53 12.66 ;
      LAYER Metal6 ;
        RECT 327.87 12 328.53 12.66 ;
      LAYER Metal3 ;
        RECT 327.87 12 328.53 12.66 ;
      LAYER Metal4 ;
        RECT 327.87 12 328.53 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 341.11 12 341.77 12.66 ;
      LAYER Metal6 ;
        RECT 341.11 12 341.77 12.66 ;
      LAYER Metal3 ;
        RECT 341.11 12 341.77 12.66 ;
      LAYER Metal4 ;
        RECT 341.11 12 341.77 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 399.1 12 399.76 12.66 ;
      LAYER Metal6 ;
        RECT 399.1 12 399.76 12.66 ;
      LAYER Metal3 ;
        RECT 399.1 12 399.76 12.66 ;
      LAYER Metal4 ;
        RECT 399.1 12 399.76 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 412.34 12 413 12.66 ;
      LAYER Metal6 ;
        RECT 412.34 12 413 12.66 ;
      LAYER Metal3 ;
        RECT 412.34 12 413 12.66 ;
      LAYER Metal4 ;
        RECT 412.34 12 413 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 441.66 12 442.32 12.66 ;
      LAYER Metal6 ;
        RECT 441.66 12 442.32 12.66 ;
      LAYER Metal3 ;
        RECT 441.66 12 442.32 12.66 ;
      LAYER Metal4 ;
        RECT 441.66 12 442.32 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 454.9 12 455.56 12.66 ;
      LAYER Metal6 ;
        RECT 454.9 12 455.56 12.66 ;
      LAYER Metal3 ;
        RECT 454.9 12 455.56 12.66 ;
      LAYER Metal4 ;
        RECT 454.9 12 455.56 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.19 12 43.85 12.66 ;
      LAYER Metal6 ;
        RECT 43.19 12 43.85 12.66 ;
      LAYER Metal3 ;
        RECT 43.19 12 43.85 12.66 ;
      LAYER Metal4 ;
        RECT 43.19 12 43.85 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 484.22 12 484.88 12.66 ;
      LAYER Metal6 ;
        RECT 484.22 12 484.88 12.66 ;
      LAYER Metal3 ;
        RECT 484.22 12 484.88 12.66 ;
      LAYER Metal4 ;
        RECT 484.22 12 484.88 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 497.46 12 498.12 12.66 ;
      LAYER Metal6 ;
        RECT 497.46 12 498.12 12.66 ;
      LAYER Metal3 ;
        RECT 497.46 12 498.12 12.66 ;
      LAYER Metal4 ;
        RECT 497.46 12 498.12 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 526.78 12 527.44 12.66 ;
      LAYER Metal6 ;
        RECT 526.78 12 527.44 12.66 ;
      LAYER Metal3 ;
        RECT 526.78 12 527.44 12.66 ;
      LAYER Metal4 ;
        RECT 526.78 12 527.44 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 540.02 12 540.68 12.66 ;
      LAYER Metal6 ;
        RECT 540.02 12 540.68 12.66 ;
      LAYER Metal3 ;
        RECT 540.02 12 540.68 12.66 ;
      LAYER Metal4 ;
        RECT 540.02 12 540.68 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 569.34 12 570 12.66 ;
      LAYER Metal6 ;
        RECT 569.34 12 570 12.66 ;
      LAYER Metal3 ;
        RECT 569.34 12 570 12.66 ;
      LAYER Metal4 ;
        RECT 569.34 12 570 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 582.58 12 583.24 12.66 ;
      LAYER Metal6 ;
        RECT 582.58 12 583.24 12.66 ;
      LAYER Metal3 ;
        RECT 582.58 12 583.24 12.66 ;
      LAYER Metal4 ;
        RECT 582.58 12 583.24 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 611.9 12 612.56 12.66 ;
      LAYER Metal6 ;
        RECT 611.9 12 612.56 12.66 ;
      LAYER Metal3 ;
        RECT 611.9 12 612.56 12.66 ;
      LAYER Metal4 ;
        RECT 611.9 12 612.56 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 625.14 12 625.8 12.66 ;
      LAYER Metal6 ;
        RECT 625.14 12 625.8 12.66 ;
      LAYER Metal3 ;
        RECT 625.14 12 625.8 12.66 ;
      LAYER Metal4 ;
        RECT 625.14 12 625.8 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 654.46 12 655.12 12.66 ;
      LAYER Metal6 ;
        RECT 654.46 12 655.12 12.66 ;
      LAYER Metal3 ;
        RECT 654.46 12 655.12 12.66 ;
      LAYER Metal4 ;
        RECT 654.46 12 655.12 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 667.7 12 668.36 12.66 ;
      LAYER Metal6 ;
        RECT 667.7 12 668.36 12.66 ;
      LAYER Metal3 ;
        RECT 667.7 12 668.36 12.66 ;
      LAYER Metal4 ;
        RECT 667.7 12 668.36 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.51 12 73.17 12.66 ;
      LAYER Metal6 ;
        RECT 72.51 12 73.17 12.66 ;
      LAYER Metal3 ;
        RECT 72.51 12 73.17 12.66 ;
      LAYER Metal4 ;
        RECT 72.51 12 73.17 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 697.02 12 697.68 12.66 ;
      LAYER Metal6 ;
        RECT 697.02 12 697.68 12.66 ;
      LAYER Metal3 ;
        RECT 697.02 12 697.68 12.66 ;
      LAYER Metal4 ;
        RECT 697.02 12 697.68 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 710.26 12 710.92 12.66 ;
      LAYER Metal6 ;
        RECT 710.26 12 710.92 12.66 ;
      LAYER Metal3 ;
        RECT 710.26 12 710.92 12.66 ;
      LAYER Metal4 ;
        RECT 710.26 12 710.92 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.75 12 86.41 12.66 ;
      LAYER Metal6 ;
        RECT 85.75 12 86.41 12.66 ;
      LAYER Metal3 ;
        RECT 85.75 12 86.41 12.66 ;
      LAYER Metal4 ;
        RECT 85.75 12 86.41 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.07 12 115.73 12.66 ;
      LAYER Metal6 ;
        RECT 115.07 12 115.73 12.66 ;
      LAYER Metal3 ;
        RECT 115.07 12 115.73 12.66 ;
      LAYER Metal4 ;
        RECT 115.07 12 115.73 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.31 12 128.97 12.66 ;
      LAYER Metal6 ;
        RECT 128.31 12 128.97 12.66 ;
      LAYER Metal3 ;
        RECT 128.31 12 128.97 12.66 ;
      LAYER Metal4 ;
        RECT 128.31 12 128.97 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.63 12 158.29 12.66 ;
      LAYER Metal6 ;
        RECT 157.63 12 158.29 12.66 ;
      LAYER Metal3 ;
        RECT 157.63 12 158.29 12.66 ;
      LAYER Metal4 ;
        RECT 157.63 12 158.29 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 170.87 12 171.53 12.66 ;
      LAYER Metal6 ;
        RECT 170.87 12 171.53 12.66 ;
      LAYER Metal3 ;
        RECT 170.87 12 171.53 12.66 ;
      LAYER Metal4 ;
        RECT 170.87 12 171.53 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 200.19 12 200.85 12.66 ;
      LAYER Metal6 ;
        RECT 200.19 12 200.85 12.66 ;
      LAYER Metal3 ;
        RECT 200.19 12 200.85 12.66 ;
      LAYER Metal4 ;
        RECT 200.19 12 200.85 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 213.43 12 214.09 12.66 ;
      LAYER Metal6 ;
        RECT 213.43 12 214.09 12.66 ;
      LAYER Metal3 ;
        RECT 213.43 12 214.09 12.66 ;
      LAYER Metal4 ;
        RECT 213.43 12 214.09 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 24.49 12 25.15 12.66 ;
      LAYER Metal6 ;
        RECT 24.49 12 25.15 12.66 ;
      LAYER Metal3 ;
        RECT 24.49 12 25.15 12.66 ;
      LAYER Metal4 ;
        RECT 24.49 12 25.15 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 237.29 12 237.95 12.66 ;
      LAYER Metal6 ;
        RECT 237.29 12 237.95 12.66 ;
      LAYER Metal3 ;
        RECT 237.29 12 237.95 12.66 ;
      LAYER Metal4 ;
        RECT 237.29 12 237.95 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 261.45 12 262.11 12.66 ;
      LAYER Metal6 ;
        RECT 261.45 12 262.11 12.66 ;
      LAYER Metal3 ;
        RECT 261.45 12 262.11 12.66 ;
      LAYER Metal4 ;
        RECT 261.45 12 262.11 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 279.85 12 280.51 12.66 ;
      LAYER Metal6 ;
        RECT 279.85 12 280.51 12.66 ;
      LAYER Metal3 ;
        RECT 279.85 12 280.51 12.66 ;
      LAYER Metal4 ;
        RECT 279.85 12 280.51 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 304.01 12 304.67 12.66 ;
      LAYER Metal6 ;
        RECT 304.01 12 304.67 12.66 ;
      LAYER Metal3 ;
        RECT 304.01 12 304.67 12.66 ;
      LAYER Metal4 ;
        RECT 304.01 12 304.67 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 322.41 12 323.07 12.66 ;
      LAYER Metal6 ;
        RECT 322.41 12 323.07 12.66 ;
      LAYER Metal3 ;
        RECT 322.41 12 323.07 12.66 ;
      LAYER Metal4 ;
        RECT 322.41 12 323.07 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 346.57 12 347.23 12.66 ;
      LAYER Metal6 ;
        RECT 346.57 12 347.23 12.66 ;
      LAYER Metal3 ;
        RECT 346.57 12 347.23 12.66 ;
      LAYER Metal4 ;
        RECT 346.57 12 347.23 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 393.64 12 394.3 12.66 ;
      LAYER Metal6 ;
        RECT 393.64 12 394.3 12.66 ;
      LAYER Metal3 ;
        RECT 393.64 12 394.3 12.66 ;
      LAYER Metal4 ;
        RECT 393.64 12 394.3 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 417.8 12 418.46 12.66 ;
      LAYER Metal6 ;
        RECT 417.8 12 418.46 12.66 ;
      LAYER Metal3 ;
        RECT 417.8 12 418.46 12.66 ;
      LAYER Metal4 ;
        RECT 417.8 12 418.46 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 436.2 12 436.86 12.66 ;
      LAYER Metal6 ;
        RECT 436.2 12 436.86 12.66 ;
      LAYER Metal3 ;
        RECT 436.2 12 436.86 12.66 ;
      LAYER Metal4 ;
        RECT 436.2 12 436.86 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 460.36 12 461.02 12.66 ;
      LAYER Metal6 ;
        RECT 460.36 12 461.02 12.66 ;
      LAYER Metal3 ;
        RECT 460.36 12 461.02 12.66 ;
      LAYER Metal4 ;
        RECT 460.36 12 461.02 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 48.65 12 49.31 12.66 ;
      LAYER Metal6 ;
        RECT 48.65 12 49.31 12.66 ;
      LAYER Metal3 ;
        RECT 48.65 12 49.31 12.66 ;
      LAYER Metal4 ;
        RECT 48.65 12 49.31 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 478.76 12 479.42 12.66 ;
      LAYER Metal6 ;
        RECT 478.76 12 479.42 12.66 ;
      LAYER Metal3 ;
        RECT 478.76 12 479.42 12.66 ;
      LAYER Metal4 ;
        RECT 478.76 12 479.42 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 502.92 12 503.58 12.66 ;
      LAYER Metal6 ;
        RECT 502.92 12 503.58 12.66 ;
      LAYER Metal3 ;
        RECT 502.92 12 503.58 12.66 ;
      LAYER Metal4 ;
        RECT 502.92 12 503.58 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 521.32 12 521.98 12.66 ;
      LAYER Metal6 ;
        RECT 521.32 12 521.98 12.66 ;
      LAYER Metal3 ;
        RECT 521.32 12 521.98 12.66 ;
      LAYER Metal4 ;
        RECT 521.32 12 521.98 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 545.48 12 546.14 12.66 ;
      LAYER Metal6 ;
        RECT 545.48 12 546.14 12.66 ;
      LAYER Metal3 ;
        RECT 545.48 12 546.14 12.66 ;
      LAYER Metal4 ;
        RECT 545.48 12 546.14 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 563.88 12 564.54 12.66 ;
      LAYER Metal6 ;
        RECT 563.88 12 564.54 12.66 ;
      LAYER Metal3 ;
        RECT 563.88 12 564.54 12.66 ;
      LAYER Metal4 ;
        RECT 563.88 12 564.54 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 588.04 12 588.7 12.66 ;
      LAYER Metal6 ;
        RECT 588.04 12 588.7 12.66 ;
      LAYER Metal3 ;
        RECT 588.04 12 588.7 12.66 ;
      LAYER Metal4 ;
        RECT 588.04 12 588.7 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 606.44 12 607.1 12.66 ;
      LAYER Metal6 ;
        RECT 606.44 12 607.1 12.66 ;
      LAYER Metal3 ;
        RECT 606.44 12 607.1 12.66 ;
      LAYER Metal4 ;
        RECT 606.44 12 607.1 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 630.6 12 631.26 12.66 ;
      LAYER Metal6 ;
        RECT 630.6 12 631.26 12.66 ;
      LAYER Metal3 ;
        RECT 630.6 12 631.26 12.66 ;
      LAYER Metal4 ;
        RECT 630.6 12 631.26 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 649 12 649.66 12.66 ;
      LAYER Metal6 ;
        RECT 649 12 649.66 12.66 ;
      LAYER Metal3 ;
        RECT 649 12 649.66 12.66 ;
      LAYER Metal4 ;
        RECT 649 12 649.66 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 673.16 12 673.82 12.66 ;
      LAYER Metal6 ;
        RECT 673.16 12 673.82 12.66 ;
      LAYER Metal3 ;
        RECT 673.16 12 673.82 12.66 ;
      LAYER Metal4 ;
        RECT 673.16 12 673.82 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.05 12 67.71 12.66 ;
      LAYER Metal6 ;
        RECT 67.05 12 67.71 12.66 ;
      LAYER Metal3 ;
        RECT 67.05 12 67.71 12.66 ;
      LAYER Metal4 ;
        RECT 67.05 12 67.71 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 691.56 12 692.22 12.66 ;
      LAYER Metal6 ;
        RECT 691.56 12 692.22 12.66 ;
      LAYER Metal3 ;
        RECT 691.56 12 692.22 12.66 ;
      LAYER Metal4 ;
        RECT 691.56 12 692.22 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 715.72 12 716.38 12.66 ;
      LAYER Metal6 ;
        RECT 715.72 12 716.38 12.66 ;
      LAYER Metal3 ;
        RECT 715.72 12 716.38 12.66 ;
      LAYER Metal4 ;
        RECT 715.72 12 716.38 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 91.21 12 91.87 12.66 ;
      LAYER Metal6 ;
        RECT 91.21 12 91.87 12.66 ;
      LAYER Metal3 ;
        RECT 91.21 12 91.87 12.66 ;
      LAYER Metal4 ;
        RECT 91.21 12 91.87 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 109.61 12 110.27 12.66 ;
      LAYER Metal6 ;
        RECT 109.61 12 110.27 12.66 ;
      LAYER Metal3 ;
        RECT 109.61 12 110.27 12.66 ;
      LAYER Metal4 ;
        RECT 109.61 12 110.27 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 133.77 12 134.43 12.66 ;
      LAYER Metal6 ;
        RECT 133.77 12 134.43 12.66 ;
      LAYER Metal3 ;
        RECT 133.77 12 134.43 12.66 ;
      LAYER Metal4 ;
        RECT 133.77 12 134.43 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 152.17 12 152.83 12.66 ;
      LAYER Metal6 ;
        RECT 152.17 12 152.83 12.66 ;
      LAYER Metal3 ;
        RECT 152.17 12 152.83 12.66 ;
      LAYER Metal4 ;
        RECT 152.17 12 152.83 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 176.33 12 176.99 12.66 ;
      LAYER Metal6 ;
        RECT 176.33 12 176.99 12.66 ;
      LAYER Metal3 ;
        RECT 176.33 12 176.99 12.66 ;
      LAYER Metal4 ;
        RECT 176.33 12 176.99 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 194.73 12 195.39 12.66 ;
      LAYER Metal6 ;
        RECT 194.73 12 195.39 12.66 ;
      LAYER Metal3 ;
        RECT 194.73 12 195.39 12.66 ;
      LAYER Metal4 ;
        RECT 194.73 12 195.39 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.89 12 219.55 12.66 ;
      LAYER Metal6 ;
        RECT 218.89 12 219.55 12.66 ;
      LAYER Metal3 ;
        RECT 218.89 12 219.55 12.66 ;
      LAYER Metal4 ;
        RECT 218.89 12 219.55 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 27.37 12 28.03 12.66 ;
      LAYER Metal6 ;
        RECT 27.37 12 28.03 12.66 ;
      LAYER Metal3 ;
        RECT 27.37 12 28.03 12.66 ;
      LAYER Metal4 ;
        RECT 27.37 12 28.03 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 240.17 12 240.83 12.66 ;
      LAYER Metal6 ;
        RECT 240.17 12 240.83 12.66 ;
      LAYER Metal3 ;
        RECT 240.17 12 240.83 12.66 ;
      LAYER Metal4 ;
        RECT 240.17 12 240.83 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 258.57 12 259.23 12.66 ;
      LAYER Metal6 ;
        RECT 258.57 12 259.23 12.66 ;
      LAYER Metal3 ;
        RECT 258.57 12 259.23 12.66 ;
      LAYER Metal4 ;
        RECT 258.57 12 259.23 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 282.73 12 283.39 12.66 ;
      LAYER Metal6 ;
        RECT 282.73 12 283.39 12.66 ;
      LAYER Metal3 ;
        RECT 282.73 12 283.39 12.66 ;
      LAYER Metal4 ;
        RECT 282.73 12 283.39 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 301.13 12 301.79 12.66 ;
      LAYER Metal6 ;
        RECT 301.13 12 301.79 12.66 ;
      LAYER Metal3 ;
        RECT 301.13 12 301.79 12.66 ;
      LAYER Metal4 ;
        RECT 301.13 12 301.79 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 325.29 12 325.95 12.66 ;
      LAYER Metal6 ;
        RECT 325.29 12 325.95 12.66 ;
      LAYER Metal3 ;
        RECT 325.29 12 325.95 12.66 ;
      LAYER Metal4 ;
        RECT 325.29 12 325.95 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 343.69 12 344.35 12.66 ;
      LAYER Metal6 ;
        RECT 343.69 12 344.35 12.66 ;
      LAYER Metal3 ;
        RECT 343.69 12 344.35 12.66 ;
      LAYER Metal4 ;
        RECT 343.69 12 344.35 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 396.52 12 397.18 12.66 ;
      LAYER Metal6 ;
        RECT 396.52 12 397.18 12.66 ;
      LAYER Metal3 ;
        RECT 396.52 12 397.18 12.66 ;
      LAYER Metal4 ;
        RECT 396.52 12 397.18 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 414.92 12 415.58 12.66 ;
      LAYER Metal6 ;
        RECT 414.92 12 415.58 12.66 ;
      LAYER Metal3 ;
        RECT 414.92 12 415.58 12.66 ;
      LAYER Metal4 ;
        RECT 414.92 12 415.58 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 439.08 12 439.74 12.66 ;
      LAYER Metal6 ;
        RECT 439.08 12 439.74 12.66 ;
      LAYER Metal3 ;
        RECT 439.08 12 439.74 12.66 ;
      LAYER Metal4 ;
        RECT 439.08 12 439.74 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 457.48 12 458.14 12.66 ;
      LAYER Metal6 ;
        RECT 457.48 12 458.14 12.66 ;
      LAYER Metal3 ;
        RECT 457.48 12 458.14 12.66 ;
      LAYER Metal4 ;
        RECT 457.48 12 458.14 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 45.77 12 46.43 12.66 ;
      LAYER Metal6 ;
        RECT 45.77 12 46.43 12.66 ;
      LAYER Metal3 ;
        RECT 45.77 12 46.43 12.66 ;
      LAYER Metal4 ;
        RECT 45.77 12 46.43 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 481.64 12 482.3 12.66 ;
      LAYER Metal6 ;
        RECT 481.64 12 482.3 12.66 ;
      LAYER Metal3 ;
        RECT 481.64 12 482.3 12.66 ;
      LAYER Metal4 ;
        RECT 481.64 12 482.3 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 500.04 12 500.7 12.66 ;
      LAYER Metal6 ;
        RECT 500.04 12 500.7 12.66 ;
      LAYER Metal3 ;
        RECT 500.04 12 500.7 12.66 ;
      LAYER Metal4 ;
        RECT 500.04 12 500.7 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 524.2 12 524.86 12.66 ;
      LAYER Metal6 ;
        RECT 524.2 12 524.86 12.66 ;
      LAYER Metal3 ;
        RECT 524.2 12 524.86 12.66 ;
      LAYER Metal4 ;
        RECT 524.2 12 524.86 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 542.6 12 543.26 12.66 ;
      LAYER Metal6 ;
        RECT 542.6 12 543.26 12.66 ;
      LAYER Metal3 ;
        RECT 542.6 12 543.26 12.66 ;
      LAYER Metal4 ;
        RECT 542.6 12 543.26 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 566.76 12 567.42 12.66 ;
      LAYER Metal6 ;
        RECT 566.76 12 567.42 12.66 ;
      LAYER Metal3 ;
        RECT 566.76 12 567.42 12.66 ;
      LAYER Metal4 ;
        RECT 566.76 12 567.42 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 585.16 12 585.82 12.66 ;
      LAYER Metal6 ;
        RECT 585.16 12 585.82 12.66 ;
      LAYER Metal3 ;
        RECT 585.16 12 585.82 12.66 ;
      LAYER Metal4 ;
        RECT 585.16 12 585.82 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 609.32 12 609.98 12.66 ;
      LAYER Metal6 ;
        RECT 609.32 12 609.98 12.66 ;
      LAYER Metal3 ;
        RECT 609.32 12 609.98 12.66 ;
      LAYER Metal4 ;
        RECT 609.32 12 609.98 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 627.72 12 628.38 12.66 ;
      LAYER Metal6 ;
        RECT 627.72 12 628.38 12.66 ;
      LAYER Metal3 ;
        RECT 627.72 12 628.38 12.66 ;
      LAYER Metal4 ;
        RECT 627.72 12 628.38 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 651.88 12 652.54 12.66 ;
      LAYER Metal6 ;
        RECT 651.88 12 652.54 12.66 ;
      LAYER Metal3 ;
        RECT 651.88 12 652.54 12.66 ;
      LAYER Metal4 ;
        RECT 651.88 12 652.54 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 670.28 12 670.94 12.66 ;
      LAYER Metal6 ;
        RECT 670.28 12 670.94 12.66 ;
      LAYER Metal3 ;
        RECT 670.28 12 670.94 12.66 ;
      LAYER Metal4 ;
        RECT 670.28 12 670.94 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.93 12 70.59 12.66 ;
      LAYER Metal6 ;
        RECT 69.93 12 70.59 12.66 ;
      LAYER Metal3 ;
        RECT 69.93 12 70.59 12.66 ;
      LAYER Metal4 ;
        RECT 69.93 12 70.59 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 694.44 12 695.1 12.66 ;
      LAYER Metal6 ;
        RECT 694.44 12 695.1 12.66 ;
      LAYER Metal3 ;
        RECT 694.44 12 695.1 12.66 ;
      LAYER Metal4 ;
        RECT 694.44 12 695.1 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 712.84 12 713.5 12.66 ;
      LAYER Metal6 ;
        RECT 712.84 12 713.5 12.66 ;
      LAYER Metal3 ;
        RECT 712.84 12 713.5 12.66 ;
      LAYER Metal4 ;
        RECT 712.84 12 713.5 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 88.33 12 88.99 12.66 ;
      LAYER Metal6 ;
        RECT 88.33 12 88.99 12.66 ;
      LAYER Metal3 ;
        RECT 88.33 12 88.99 12.66 ;
      LAYER Metal4 ;
        RECT 88.33 12 88.99 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 112.49 12 113.15 12.66 ;
      LAYER Metal6 ;
        RECT 112.49 12 113.15 12.66 ;
      LAYER Metal3 ;
        RECT 112.49 12 113.15 12.66 ;
      LAYER Metal4 ;
        RECT 112.49 12 113.15 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 130.89 12 131.55 12.66 ;
      LAYER Metal6 ;
        RECT 130.89 12 131.55 12.66 ;
      LAYER Metal3 ;
        RECT 130.89 12 131.55 12.66 ;
      LAYER Metal4 ;
        RECT 130.89 12 131.55 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 155.05 12 155.71 12.66 ;
      LAYER Metal6 ;
        RECT 155.05 12 155.71 12.66 ;
      LAYER Metal3 ;
        RECT 155.05 12 155.71 12.66 ;
      LAYER Metal4 ;
        RECT 155.05 12 155.71 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 173.45 12 174.11 12.66 ;
      LAYER Metal6 ;
        RECT 173.45 12 174.11 12.66 ;
      LAYER Metal3 ;
        RECT 173.45 12 174.11 12.66 ;
      LAYER Metal4 ;
        RECT 173.45 12 174.11 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 197.61 12 198.27 12.66 ;
      LAYER Metal6 ;
        RECT 197.61 12 198.27 12.66 ;
      LAYER Metal3 ;
        RECT 197.61 12 198.27 12.66 ;
      LAYER Metal4 ;
        RECT 197.61 12 198.27 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 216.01 12 216.67 12.66 ;
      LAYER Metal6 ;
        RECT 216.01 12 216.67 12.66 ;
      LAYER Metal3 ;
        RECT 216.01 12 216.67 12.66 ;
      LAYER Metal4 ;
        RECT 216.01 12 216.67 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.01 12 376.67 12.66 ;
      LAYER Metal6 ;
        RECT 376.01 12 376.67 12.66 ;
      LAYER Metal3 ;
        RECT 376.01 12 376.67 12.66 ;
      LAYER Metal4 ;
        RECT 376.01 12 376.67 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 364.2 12 364.86 12.66 ;
      LAYER Metal6 ;
        RECT 364.2 12 364.86 12.66 ;
      LAYER Metal3 ;
        RECT 364.2 12 364.86 12.66 ;
      LAYER Metal4 ;
        RECT 364.2 12 364.86 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 517.75 761.745 522.75 ;
        RECT 0 0 761.745 5 ;
      LAYER Metal2 ;
        RECT 756.745 0 761.745 522.75 ;
        RECT 0 0 5 522.75 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 512.15 756.145 517.15 ;
        RECT 5.6 5.6 756.145 10.6 ;
      LAYER Metal2 ;
        RECT 751.145 5.6 756.145 517.15 ;
        RECT 5.6 5.6 10.6 517.15 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 749.79 510.725 ;
    LAYER Metal2 ;
      RECT 12 12 749.79 510.725 ;
    LAYER Metal3 ;
      RECT 12 12 749.79 510.725 ;
    LAYER Metal4 ;
      RECT 12 12 749.79 510.725 ;
    LAYER Metal5 ;
      RECT 12 12 749.79 510.725 ;
    LAYER Metal6 ;
      RECT 12 12 749.79 510.725 ;
  END
END MEM2_2048X32

END LIBRARY
