VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MEM2_1024X32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2_1024X32 0 0 ;
  SIZE 772.885 BY 307.3 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 216.54 12.66 217.2 ;
      LAYER Metal6 ;
        RECT 12 216.54 12.66 217.2 ;
      LAYER Metal3 ;
        RECT 12 216.54 12.66 217.2 ;
      LAYER Metal4 ;
        RECT 12 216.54 12.66 217.2 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 210.42 12.66 211.08 ;
      LAYER Metal6 ;
        RECT 12 210.42 12.66 211.08 ;
      LAYER Metal3 ;
        RECT 12 210.42 12.66 211.08 ;
      LAYER Metal4 ;
        RECT 12 210.42 12.66 211.08 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 207.32 12.66 207.98 ;
      LAYER Metal6 ;
        RECT 12 207.32 12.66 207.98 ;
      LAYER Metal3 ;
        RECT 12 207.32 12.66 207.98 ;
      LAYER Metal4 ;
        RECT 12 207.32 12.66 207.98 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 201.2 12.66 201.86 ;
      LAYER Metal6 ;
        RECT 12 201.2 12.66 201.86 ;
      LAYER Metal3 ;
        RECT 12 201.2 12.66 201.86 ;
      LAYER Metal4 ;
        RECT 12 201.2 12.66 201.86 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 198.18 12.66 198.84 ;
      LAYER Metal6 ;
        RECT 12 198.18 12.66 198.84 ;
      LAYER Metal3 ;
        RECT 12 198.18 12.66 198.84 ;
      LAYER Metal4 ;
        RECT 12 198.18 12.66 198.84 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 195.08 12.66 195.74 ;
      LAYER Metal6 ;
        RECT 12 195.08 12.66 195.74 ;
      LAYER Metal3 ;
        RECT 12 195.08 12.66 195.74 ;
      LAYER Metal4 ;
        RECT 12 195.08 12.66 195.74 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 188.96 12.66 189.62 ;
      LAYER Metal6 ;
        RECT 12 188.96 12.66 189.62 ;
      LAYER Metal3 ;
        RECT 12 188.96 12.66 189.62 ;
      LAYER Metal4 ;
        RECT 12 188.96 12.66 189.62 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 185.94 12.66 186.6 ;
      LAYER Metal6 ;
        RECT 12 185.94 12.66 186.6 ;
      LAYER Metal3 ;
        RECT 12 185.94 12.66 186.6 ;
      LAYER Metal4 ;
        RECT 12 185.94 12.66 186.6 ;
    END
  END A1[7]
  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 182.84 12.66 183.5 ;
      LAYER Metal6 ;
        RECT 12 182.84 12.66 183.5 ;
      LAYER Metal3 ;
        RECT 12 182.84 12.66 183.5 ;
      LAYER Metal4 ;
        RECT 12 182.84 12.66 183.5 ;
    END
  END A1[8]
  PIN A1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 176.72 12.66 177.38 ;
      LAYER Metal6 ;
        RECT 12 176.72 12.66 177.38 ;
      LAYER Metal3 ;
        RECT 12 176.72 12.66 177.38 ;
      LAYER Metal4 ;
        RECT 12 176.72 12.66 177.38 ;
    END
  END A1[9]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 132.16 12.66 132.82 ;
      LAYER Metal6 ;
        RECT 12 132.16 12.66 132.82 ;
      LAYER Metal3 ;
        RECT 12 132.16 12.66 132.82 ;
      LAYER Metal4 ;
        RECT 12 132.16 12.66 132.82 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 138.28 12.66 138.94 ;
      LAYER Metal6 ;
        RECT 12 138.28 12.66 138.94 ;
      LAYER Metal3 ;
        RECT 12 138.28 12.66 138.94 ;
      LAYER Metal4 ;
        RECT 12 138.28 12.66 138.94 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 141.38 12.66 142.04 ;
      LAYER Metal6 ;
        RECT 12 141.38 12.66 142.04 ;
      LAYER Metal3 ;
        RECT 12 141.38 12.66 142.04 ;
      LAYER Metal4 ;
        RECT 12 141.38 12.66 142.04 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 147.5 12.66 148.16 ;
      LAYER Metal6 ;
        RECT 12 147.5 12.66 148.16 ;
      LAYER Metal3 ;
        RECT 12 147.5 12.66 148.16 ;
      LAYER Metal4 ;
        RECT 12 147.5 12.66 148.16 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 150.52 12.66 151.18 ;
      LAYER Metal6 ;
        RECT 12 150.52 12.66 151.18 ;
      LAYER Metal3 ;
        RECT 12 150.52 12.66 151.18 ;
      LAYER Metal4 ;
        RECT 12 150.52 12.66 151.18 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 153.62 12.66 154.28 ;
      LAYER Metal6 ;
        RECT 12 153.62 12.66 154.28 ;
      LAYER Metal3 ;
        RECT 12 153.62 12.66 154.28 ;
      LAYER Metal4 ;
        RECT 12 153.62 12.66 154.28 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 159.74 12.66 160.4 ;
      LAYER Metal6 ;
        RECT 12 159.74 12.66 160.4 ;
      LAYER Metal3 ;
        RECT 12 159.74 12.66 160.4 ;
      LAYER Metal4 ;
        RECT 12 159.74 12.66 160.4 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 162.76 12.66 163.42 ;
      LAYER Metal6 ;
        RECT 12 162.76 12.66 163.42 ;
      LAYER Metal3 ;
        RECT 12 162.76 12.66 163.42 ;
      LAYER Metal4 ;
        RECT 12 162.76 12.66 163.42 ;
    END
  END A2[7]
  PIN A2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 165.86 12.66 166.52 ;
      LAYER Metal6 ;
        RECT 12 165.86 12.66 166.52 ;
      LAYER Metal3 ;
        RECT 12 165.86 12.66 166.52 ;
      LAYER Metal4 ;
        RECT 12 165.86 12.66 166.52 ;
    END
  END A2[8]
  PIN A2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 171.98 12.66 172.64 ;
      LAYER Metal6 ;
        RECT 12 171.98 12.66 172.64 ;
      LAYER Metal3 ;
        RECT 12 171.98 12.66 172.64 ;
      LAYER Metal4 ;
        RECT 12 171.98 12.66 172.64 ;
    END
  END A2[9]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 382.025 12 382.685 12.66 ;
      LAYER Metal6 ;
        RECT 382.025 12 382.685 12.66 ;
      LAYER Metal3 ;
        RECT 382.025 12 382.685 12.66 ;
      LAYER Metal4 ;
        RECT 382.025 12 382.685 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.6 12 367.26 12.66 ;
      LAYER Metal6 ;
        RECT 366.6 12 367.26 12.66 ;
      LAYER Metal3 ;
        RECT 366.6 12 367.26 12.66 ;
      LAYER Metal4 ;
        RECT 366.6 12 367.26 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 390.65 12 391.31 12.66 ;
      LAYER Metal6 ;
        RECT 390.65 12 391.31 12.66 ;
      LAYER Metal3 ;
        RECT 390.65 12 391.31 12.66 ;
      LAYER Metal4 ;
        RECT 390.65 12 391.31 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 357.975 12 358.635 12.66 ;
      LAYER Metal6 ;
        RECT 357.975 12 358.635 12.66 ;
      LAYER Metal3 ;
        RECT 357.975 12 358.635 12.66 ;
      LAYER Metal4 ;
        RECT 357.975 12 358.635 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 21.91 12 22.57 12.66 ;
      LAYER Metal6 ;
        RECT 21.91 12 22.57 12.66 ;
      LAYER Metal3 ;
        RECT 21.91 12 22.57 12.66 ;
      LAYER Metal4 ;
        RECT 21.91 12 22.57 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 234.71 12 235.37 12.66 ;
      LAYER Metal6 ;
        RECT 234.71 12 235.37 12.66 ;
      LAYER Metal3 ;
        RECT 234.71 12 235.37 12.66 ;
      LAYER Metal4 ;
        RECT 234.71 12 235.37 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.03 12 264.69 12.66 ;
      LAYER Metal6 ;
        RECT 264.03 12 264.69 12.66 ;
      LAYER Metal3 ;
        RECT 264.03 12 264.69 12.66 ;
      LAYER Metal4 ;
        RECT 264.03 12 264.69 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 277.27 12 277.93 12.66 ;
      LAYER Metal6 ;
        RECT 277.27 12 277.93 12.66 ;
      LAYER Metal3 ;
        RECT 277.27 12 277.93 12.66 ;
      LAYER Metal4 ;
        RECT 277.27 12 277.93 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.59 12 307.25 12.66 ;
      LAYER Metal6 ;
        RECT 306.59 12 307.25 12.66 ;
      LAYER Metal3 ;
        RECT 306.59 12 307.25 12.66 ;
      LAYER Metal4 ;
        RECT 306.59 12 307.25 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 319.83 12 320.49 12.66 ;
      LAYER Metal6 ;
        RECT 319.83 12 320.49 12.66 ;
      LAYER Metal3 ;
        RECT 319.83 12 320.49 12.66 ;
      LAYER Metal4 ;
        RECT 319.83 12 320.49 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.15 12 349.81 12.66 ;
      LAYER Metal6 ;
        RECT 349.15 12 349.81 12.66 ;
      LAYER Metal3 ;
        RECT 349.15 12 349.81 12.66 ;
      LAYER Metal4 ;
        RECT 349.15 12 349.81 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 399.475 12 400.135 12.66 ;
      LAYER Metal6 ;
        RECT 399.475 12 400.135 12.66 ;
      LAYER Metal3 ;
        RECT 399.475 12 400.135 12.66 ;
      LAYER Metal4 ;
        RECT 399.475 12 400.135 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 428.795 12 429.455 12.66 ;
      LAYER Metal6 ;
        RECT 428.795 12 429.455 12.66 ;
      LAYER Metal3 ;
        RECT 428.795 12 429.455 12.66 ;
      LAYER Metal4 ;
        RECT 428.795 12 429.455 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 442.035 12 442.695 12.66 ;
      LAYER Metal6 ;
        RECT 442.035 12 442.695 12.66 ;
      LAYER Metal3 ;
        RECT 442.035 12 442.695 12.66 ;
      LAYER Metal4 ;
        RECT 442.035 12 442.695 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 471.355 12 472.015 12.66 ;
      LAYER Metal6 ;
        RECT 471.355 12 472.015 12.66 ;
      LAYER Metal3 ;
        RECT 471.355 12 472.015 12.66 ;
      LAYER Metal4 ;
        RECT 471.355 12 472.015 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.23 12 51.89 12.66 ;
      LAYER Metal6 ;
        RECT 51.23 12 51.89 12.66 ;
      LAYER Metal3 ;
        RECT 51.23 12 51.89 12.66 ;
      LAYER Metal4 ;
        RECT 51.23 12 51.89 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 484.595 12 485.255 12.66 ;
      LAYER Metal6 ;
        RECT 484.595 12 485.255 12.66 ;
      LAYER Metal3 ;
        RECT 484.595 12 485.255 12.66 ;
      LAYER Metal4 ;
        RECT 484.595 12 485.255 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 513.915 12 514.575 12.66 ;
      LAYER Metal6 ;
        RECT 513.915 12 514.575 12.66 ;
      LAYER Metal3 ;
        RECT 513.915 12 514.575 12.66 ;
      LAYER Metal4 ;
        RECT 513.915 12 514.575 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 527.155 12 527.815 12.66 ;
      LAYER Metal6 ;
        RECT 527.155 12 527.815 12.66 ;
      LAYER Metal3 ;
        RECT 527.155 12 527.815 12.66 ;
      LAYER Metal4 ;
        RECT 527.155 12 527.815 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 556.475 12 557.135 12.66 ;
      LAYER Metal6 ;
        RECT 556.475 12 557.135 12.66 ;
      LAYER Metal3 ;
        RECT 556.475 12 557.135 12.66 ;
      LAYER Metal4 ;
        RECT 556.475 12 557.135 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 569.715 12 570.375 12.66 ;
      LAYER Metal6 ;
        RECT 569.715 12 570.375 12.66 ;
      LAYER Metal3 ;
        RECT 569.715 12 570.375 12.66 ;
      LAYER Metal4 ;
        RECT 569.715 12 570.375 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 599.035 12 599.695 12.66 ;
      LAYER Metal6 ;
        RECT 599.035 12 599.695 12.66 ;
      LAYER Metal3 ;
        RECT 599.035 12 599.695 12.66 ;
      LAYER Metal4 ;
        RECT 599.035 12 599.695 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 612.275 12 612.935 12.66 ;
      LAYER Metal6 ;
        RECT 612.275 12 612.935 12.66 ;
      LAYER Metal3 ;
        RECT 612.275 12 612.935 12.66 ;
      LAYER Metal4 ;
        RECT 612.275 12 612.935 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 641.595 12 642.255 12.66 ;
      LAYER Metal6 ;
        RECT 641.595 12 642.255 12.66 ;
      LAYER Metal3 ;
        RECT 641.595 12 642.255 12.66 ;
      LAYER Metal4 ;
        RECT 641.595 12 642.255 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 654.835 12 655.495 12.66 ;
      LAYER Metal6 ;
        RECT 654.835 12 655.495 12.66 ;
      LAYER Metal3 ;
        RECT 654.835 12 655.495 12.66 ;
      LAYER Metal4 ;
        RECT 654.835 12 655.495 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 684.155 12 684.815 12.66 ;
      LAYER Metal6 ;
        RECT 684.155 12 684.815 12.66 ;
      LAYER Metal3 ;
        RECT 684.155 12 684.815 12.66 ;
      LAYER Metal4 ;
        RECT 684.155 12 684.815 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.47 12 65.13 12.66 ;
      LAYER Metal6 ;
        RECT 64.47 12 65.13 12.66 ;
      LAYER Metal3 ;
        RECT 64.47 12 65.13 12.66 ;
      LAYER Metal4 ;
        RECT 64.47 12 65.13 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 697.395 12 698.055 12.66 ;
      LAYER Metal6 ;
        RECT 697.395 12 698.055 12.66 ;
      LAYER Metal3 ;
        RECT 697.395 12 698.055 12.66 ;
      LAYER Metal4 ;
        RECT 697.395 12 698.055 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 726.715 12 727.375 12.66 ;
      LAYER Metal6 ;
        RECT 726.715 12 727.375 12.66 ;
      LAYER Metal3 ;
        RECT 726.715 12 727.375 12.66 ;
      LAYER Metal4 ;
        RECT 726.715 12 727.375 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.79 12 94.45 12.66 ;
      LAYER Metal6 ;
        RECT 93.79 12 94.45 12.66 ;
      LAYER Metal3 ;
        RECT 93.79 12 94.45 12.66 ;
      LAYER Metal4 ;
        RECT 93.79 12 94.45 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.03 12 107.69 12.66 ;
      LAYER Metal6 ;
        RECT 107.03 12 107.69 12.66 ;
      LAYER Metal3 ;
        RECT 107.03 12 107.69 12.66 ;
      LAYER Metal4 ;
        RECT 107.03 12 107.69 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.35 12 137.01 12.66 ;
      LAYER Metal6 ;
        RECT 136.35 12 137.01 12.66 ;
      LAYER Metal3 ;
        RECT 136.35 12 137.01 12.66 ;
      LAYER Metal4 ;
        RECT 136.35 12 137.01 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.59 12 150.25 12.66 ;
      LAYER Metal6 ;
        RECT 149.59 12 150.25 12.66 ;
      LAYER Metal3 ;
        RECT 149.59 12 150.25 12.66 ;
      LAYER Metal4 ;
        RECT 149.59 12 150.25 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.91 12 179.57 12.66 ;
      LAYER Metal6 ;
        RECT 178.91 12 179.57 12.66 ;
      LAYER Metal3 ;
        RECT 178.91 12 179.57 12.66 ;
      LAYER Metal4 ;
        RECT 178.91 12 179.57 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 192.15 12 192.81 12.66 ;
      LAYER Metal6 ;
        RECT 192.15 12 192.81 12.66 ;
      LAYER Metal3 ;
        RECT 192.15 12 192.81 12.66 ;
      LAYER Metal4 ;
        RECT 192.15 12 192.81 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.47 12 222.13 12.66 ;
      LAYER Metal6 ;
        RECT 221.47 12 222.13 12.66 ;
      LAYER Metal3 ;
        RECT 221.47 12 222.13 12.66 ;
      LAYER Metal4 ;
        RECT 221.47 12 222.13 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.95 12 30.61 12.66 ;
      LAYER Metal6 ;
        RECT 29.95 12 30.61 12.66 ;
      LAYER Metal3 ;
        RECT 29.95 12 30.61 12.66 ;
      LAYER Metal4 ;
        RECT 29.95 12 30.61 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.75 12 243.41 12.66 ;
      LAYER Metal6 ;
        RECT 242.75 12 243.41 12.66 ;
      LAYER Metal3 ;
        RECT 242.75 12 243.41 12.66 ;
      LAYER Metal4 ;
        RECT 242.75 12 243.41 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 255.99 12 256.65 12.66 ;
      LAYER Metal6 ;
        RECT 255.99 12 256.65 12.66 ;
      LAYER Metal3 ;
        RECT 255.99 12 256.65 12.66 ;
      LAYER Metal4 ;
        RECT 255.99 12 256.65 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.31 12 285.97 12.66 ;
      LAYER Metal6 ;
        RECT 285.31 12 285.97 12.66 ;
      LAYER Metal3 ;
        RECT 285.31 12 285.97 12.66 ;
      LAYER Metal4 ;
        RECT 285.31 12 285.97 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 298.55 12 299.21 12.66 ;
      LAYER Metal6 ;
        RECT 298.55 12 299.21 12.66 ;
      LAYER Metal3 ;
        RECT 298.55 12 299.21 12.66 ;
      LAYER Metal4 ;
        RECT 298.55 12 299.21 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 327.87 12 328.53 12.66 ;
      LAYER Metal6 ;
        RECT 327.87 12 328.53 12.66 ;
      LAYER Metal3 ;
        RECT 327.87 12 328.53 12.66 ;
      LAYER Metal4 ;
        RECT 327.87 12 328.53 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 341.11 12 341.77 12.66 ;
      LAYER Metal6 ;
        RECT 341.11 12 341.77 12.66 ;
      LAYER Metal3 ;
        RECT 341.11 12 341.77 12.66 ;
      LAYER Metal4 ;
        RECT 341.11 12 341.77 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 407.515 12 408.175 12.66 ;
      LAYER Metal6 ;
        RECT 407.515 12 408.175 12.66 ;
      LAYER Metal3 ;
        RECT 407.515 12 408.175 12.66 ;
      LAYER Metal4 ;
        RECT 407.515 12 408.175 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 420.755 12 421.415 12.66 ;
      LAYER Metal6 ;
        RECT 420.755 12 421.415 12.66 ;
      LAYER Metal3 ;
        RECT 420.755 12 421.415 12.66 ;
      LAYER Metal4 ;
        RECT 420.755 12 421.415 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 450.075 12 450.735 12.66 ;
      LAYER Metal6 ;
        RECT 450.075 12 450.735 12.66 ;
      LAYER Metal3 ;
        RECT 450.075 12 450.735 12.66 ;
      LAYER Metal4 ;
        RECT 450.075 12 450.735 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 463.315 12 463.975 12.66 ;
      LAYER Metal6 ;
        RECT 463.315 12 463.975 12.66 ;
      LAYER Metal3 ;
        RECT 463.315 12 463.975 12.66 ;
      LAYER Metal4 ;
        RECT 463.315 12 463.975 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.19 12 43.85 12.66 ;
      LAYER Metal6 ;
        RECT 43.19 12 43.85 12.66 ;
      LAYER Metal3 ;
        RECT 43.19 12 43.85 12.66 ;
      LAYER Metal4 ;
        RECT 43.19 12 43.85 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 492.635 12 493.295 12.66 ;
      LAYER Metal6 ;
        RECT 492.635 12 493.295 12.66 ;
      LAYER Metal3 ;
        RECT 492.635 12 493.295 12.66 ;
      LAYER Metal4 ;
        RECT 492.635 12 493.295 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 505.875 12 506.535 12.66 ;
      LAYER Metal6 ;
        RECT 505.875 12 506.535 12.66 ;
      LAYER Metal3 ;
        RECT 505.875 12 506.535 12.66 ;
      LAYER Metal4 ;
        RECT 505.875 12 506.535 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 535.195 12 535.855 12.66 ;
      LAYER Metal6 ;
        RECT 535.195 12 535.855 12.66 ;
      LAYER Metal3 ;
        RECT 535.195 12 535.855 12.66 ;
      LAYER Metal4 ;
        RECT 535.195 12 535.855 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 548.435 12 549.095 12.66 ;
      LAYER Metal6 ;
        RECT 548.435 12 549.095 12.66 ;
      LAYER Metal3 ;
        RECT 548.435 12 549.095 12.66 ;
      LAYER Metal4 ;
        RECT 548.435 12 549.095 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 577.755 12 578.415 12.66 ;
      LAYER Metal6 ;
        RECT 577.755 12 578.415 12.66 ;
      LAYER Metal3 ;
        RECT 577.755 12 578.415 12.66 ;
      LAYER Metal4 ;
        RECT 577.755 12 578.415 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 590.995 12 591.655 12.66 ;
      LAYER Metal6 ;
        RECT 590.995 12 591.655 12.66 ;
      LAYER Metal3 ;
        RECT 590.995 12 591.655 12.66 ;
      LAYER Metal4 ;
        RECT 590.995 12 591.655 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 620.315 12 620.975 12.66 ;
      LAYER Metal6 ;
        RECT 620.315 12 620.975 12.66 ;
      LAYER Metal3 ;
        RECT 620.315 12 620.975 12.66 ;
      LAYER Metal4 ;
        RECT 620.315 12 620.975 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 633.555 12 634.215 12.66 ;
      LAYER Metal6 ;
        RECT 633.555 12 634.215 12.66 ;
      LAYER Metal3 ;
        RECT 633.555 12 634.215 12.66 ;
      LAYER Metal4 ;
        RECT 633.555 12 634.215 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 662.875 12 663.535 12.66 ;
      LAYER Metal6 ;
        RECT 662.875 12 663.535 12.66 ;
      LAYER Metal3 ;
        RECT 662.875 12 663.535 12.66 ;
      LAYER Metal4 ;
        RECT 662.875 12 663.535 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 676.115 12 676.775 12.66 ;
      LAYER Metal6 ;
        RECT 676.115 12 676.775 12.66 ;
      LAYER Metal3 ;
        RECT 676.115 12 676.775 12.66 ;
      LAYER Metal4 ;
        RECT 676.115 12 676.775 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.51 12 73.17 12.66 ;
      LAYER Metal6 ;
        RECT 72.51 12 73.17 12.66 ;
      LAYER Metal3 ;
        RECT 72.51 12 73.17 12.66 ;
      LAYER Metal4 ;
        RECT 72.51 12 73.17 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 705.435 12 706.095 12.66 ;
      LAYER Metal6 ;
        RECT 705.435 12 706.095 12.66 ;
      LAYER Metal3 ;
        RECT 705.435 12 706.095 12.66 ;
      LAYER Metal4 ;
        RECT 705.435 12 706.095 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 718.675 12 719.335 12.66 ;
      LAYER Metal6 ;
        RECT 718.675 12 719.335 12.66 ;
      LAYER Metal3 ;
        RECT 718.675 12 719.335 12.66 ;
      LAYER Metal4 ;
        RECT 718.675 12 719.335 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.75 12 86.41 12.66 ;
      LAYER Metal6 ;
        RECT 85.75 12 86.41 12.66 ;
      LAYER Metal3 ;
        RECT 85.75 12 86.41 12.66 ;
      LAYER Metal4 ;
        RECT 85.75 12 86.41 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.07 12 115.73 12.66 ;
      LAYER Metal6 ;
        RECT 115.07 12 115.73 12.66 ;
      LAYER Metal3 ;
        RECT 115.07 12 115.73 12.66 ;
      LAYER Metal4 ;
        RECT 115.07 12 115.73 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.31 12 128.97 12.66 ;
      LAYER Metal6 ;
        RECT 128.31 12 128.97 12.66 ;
      LAYER Metal3 ;
        RECT 128.31 12 128.97 12.66 ;
      LAYER Metal4 ;
        RECT 128.31 12 128.97 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.63 12 158.29 12.66 ;
      LAYER Metal6 ;
        RECT 157.63 12 158.29 12.66 ;
      LAYER Metal3 ;
        RECT 157.63 12 158.29 12.66 ;
      LAYER Metal4 ;
        RECT 157.63 12 158.29 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 170.87 12 171.53 12.66 ;
      LAYER Metal6 ;
        RECT 170.87 12 171.53 12.66 ;
      LAYER Metal3 ;
        RECT 170.87 12 171.53 12.66 ;
      LAYER Metal4 ;
        RECT 170.87 12 171.53 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 200.19 12 200.85 12.66 ;
      LAYER Metal6 ;
        RECT 200.19 12 200.85 12.66 ;
      LAYER Metal3 ;
        RECT 200.19 12 200.85 12.66 ;
      LAYER Metal4 ;
        RECT 200.19 12 200.85 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 213.43 12 214.09 12.66 ;
      LAYER Metal6 ;
        RECT 213.43 12 214.09 12.66 ;
      LAYER Metal3 ;
        RECT 213.43 12 214.09 12.66 ;
      LAYER Metal4 ;
        RECT 213.43 12 214.09 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 24.49 12 25.15 12.66 ;
      LAYER Metal6 ;
        RECT 24.49 12 25.15 12.66 ;
      LAYER Metal3 ;
        RECT 24.49 12 25.15 12.66 ;
      LAYER Metal4 ;
        RECT 24.49 12 25.15 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 237.29 12 237.95 12.66 ;
      LAYER Metal6 ;
        RECT 237.29 12 237.95 12.66 ;
      LAYER Metal3 ;
        RECT 237.29 12 237.95 12.66 ;
      LAYER Metal4 ;
        RECT 237.29 12 237.95 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 261.45 12 262.11 12.66 ;
      LAYER Metal6 ;
        RECT 261.45 12 262.11 12.66 ;
      LAYER Metal3 ;
        RECT 261.45 12 262.11 12.66 ;
      LAYER Metal4 ;
        RECT 261.45 12 262.11 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 279.85 12 280.51 12.66 ;
      LAYER Metal6 ;
        RECT 279.85 12 280.51 12.66 ;
      LAYER Metal3 ;
        RECT 279.85 12 280.51 12.66 ;
      LAYER Metal4 ;
        RECT 279.85 12 280.51 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 304.01 12 304.67 12.66 ;
      LAYER Metal6 ;
        RECT 304.01 12 304.67 12.66 ;
      LAYER Metal3 ;
        RECT 304.01 12 304.67 12.66 ;
      LAYER Metal4 ;
        RECT 304.01 12 304.67 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 322.41 12 323.07 12.66 ;
      LAYER Metal6 ;
        RECT 322.41 12 323.07 12.66 ;
      LAYER Metal3 ;
        RECT 322.41 12 323.07 12.66 ;
      LAYER Metal4 ;
        RECT 322.41 12 323.07 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 346.57 12 347.23 12.66 ;
      LAYER Metal6 ;
        RECT 346.57 12 347.23 12.66 ;
      LAYER Metal3 ;
        RECT 346.57 12 347.23 12.66 ;
      LAYER Metal4 ;
        RECT 346.57 12 347.23 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 402.055 12 402.715 12.66 ;
      LAYER Metal6 ;
        RECT 402.055 12 402.715 12.66 ;
      LAYER Metal3 ;
        RECT 402.055 12 402.715 12.66 ;
      LAYER Metal4 ;
        RECT 402.055 12 402.715 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 426.215 12 426.875 12.66 ;
      LAYER Metal6 ;
        RECT 426.215 12 426.875 12.66 ;
      LAYER Metal3 ;
        RECT 426.215 12 426.875 12.66 ;
      LAYER Metal4 ;
        RECT 426.215 12 426.875 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 444.615 12 445.275 12.66 ;
      LAYER Metal6 ;
        RECT 444.615 12 445.275 12.66 ;
      LAYER Metal3 ;
        RECT 444.615 12 445.275 12.66 ;
      LAYER Metal4 ;
        RECT 444.615 12 445.275 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 468.775 12 469.435 12.66 ;
      LAYER Metal6 ;
        RECT 468.775 12 469.435 12.66 ;
      LAYER Metal3 ;
        RECT 468.775 12 469.435 12.66 ;
      LAYER Metal4 ;
        RECT 468.775 12 469.435 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 48.65 12 49.31 12.66 ;
      LAYER Metal6 ;
        RECT 48.65 12 49.31 12.66 ;
      LAYER Metal3 ;
        RECT 48.65 12 49.31 12.66 ;
      LAYER Metal4 ;
        RECT 48.65 12 49.31 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 487.175 12 487.835 12.66 ;
      LAYER Metal6 ;
        RECT 487.175 12 487.835 12.66 ;
      LAYER Metal3 ;
        RECT 487.175 12 487.835 12.66 ;
      LAYER Metal4 ;
        RECT 487.175 12 487.835 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 511.335 12 511.995 12.66 ;
      LAYER Metal6 ;
        RECT 511.335 12 511.995 12.66 ;
      LAYER Metal3 ;
        RECT 511.335 12 511.995 12.66 ;
      LAYER Metal4 ;
        RECT 511.335 12 511.995 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 529.735 12 530.395 12.66 ;
      LAYER Metal6 ;
        RECT 529.735 12 530.395 12.66 ;
      LAYER Metal3 ;
        RECT 529.735 12 530.395 12.66 ;
      LAYER Metal4 ;
        RECT 529.735 12 530.395 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 553.895 12 554.555 12.66 ;
      LAYER Metal6 ;
        RECT 553.895 12 554.555 12.66 ;
      LAYER Metal3 ;
        RECT 553.895 12 554.555 12.66 ;
      LAYER Metal4 ;
        RECT 553.895 12 554.555 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 572.295 12 572.955 12.66 ;
      LAYER Metal6 ;
        RECT 572.295 12 572.955 12.66 ;
      LAYER Metal3 ;
        RECT 572.295 12 572.955 12.66 ;
      LAYER Metal4 ;
        RECT 572.295 12 572.955 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 596.455 12 597.115 12.66 ;
      LAYER Metal6 ;
        RECT 596.455 12 597.115 12.66 ;
      LAYER Metal3 ;
        RECT 596.455 12 597.115 12.66 ;
      LAYER Metal4 ;
        RECT 596.455 12 597.115 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 614.855 12 615.515 12.66 ;
      LAYER Metal6 ;
        RECT 614.855 12 615.515 12.66 ;
      LAYER Metal3 ;
        RECT 614.855 12 615.515 12.66 ;
      LAYER Metal4 ;
        RECT 614.855 12 615.515 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 639.015 12 639.675 12.66 ;
      LAYER Metal6 ;
        RECT 639.015 12 639.675 12.66 ;
      LAYER Metal3 ;
        RECT 639.015 12 639.675 12.66 ;
      LAYER Metal4 ;
        RECT 639.015 12 639.675 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 657.415 12 658.075 12.66 ;
      LAYER Metal6 ;
        RECT 657.415 12 658.075 12.66 ;
      LAYER Metal3 ;
        RECT 657.415 12 658.075 12.66 ;
      LAYER Metal4 ;
        RECT 657.415 12 658.075 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 681.575 12 682.235 12.66 ;
      LAYER Metal6 ;
        RECT 681.575 12 682.235 12.66 ;
      LAYER Metal3 ;
        RECT 681.575 12 682.235 12.66 ;
      LAYER Metal4 ;
        RECT 681.575 12 682.235 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.05 12 67.71 12.66 ;
      LAYER Metal6 ;
        RECT 67.05 12 67.71 12.66 ;
      LAYER Metal3 ;
        RECT 67.05 12 67.71 12.66 ;
      LAYER Metal4 ;
        RECT 67.05 12 67.71 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 699.975 12 700.635 12.66 ;
      LAYER Metal6 ;
        RECT 699.975 12 700.635 12.66 ;
      LAYER Metal3 ;
        RECT 699.975 12 700.635 12.66 ;
      LAYER Metal4 ;
        RECT 699.975 12 700.635 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 724.135 12 724.795 12.66 ;
      LAYER Metal6 ;
        RECT 724.135 12 724.795 12.66 ;
      LAYER Metal3 ;
        RECT 724.135 12 724.795 12.66 ;
      LAYER Metal4 ;
        RECT 724.135 12 724.795 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 91.21 12 91.87 12.66 ;
      LAYER Metal6 ;
        RECT 91.21 12 91.87 12.66 ;
      LAYER Metal3 ;
        RECT 91.21 12 91.87 12.66 ;
      LAYER Metal4 ;
        RECT 91.21 12 91.87 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 109.61 12 110.27 12.66 ;
      LAYER Metal6 ;
        RECT 109.61 12 110.27 12.66 ;
      LAYER Metal3 ;
        RECT 109.61 12 110.27 12.66 ;
      LAYER Metal4 ;
        RECT 109.61 12 110.27 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 133.77 12 134.43 12.66 ;
      LAYER Metal6 ;
        RECT 133.77 12 134.43 12.66 ;
      LAYER Metal3 ;
        RECT 133.77 12 134.43 12.66 ;
      LAYER Metal4 ;
        RECT 133.77 12 134.43 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 152.17 12 152.83 12.66 ;
      LAYER Metal6 ;
        RECT 152.17 12 152.83 12.66 ;
      LAYER Metal3 ;
        RECT 152.17 12 152.83 12.66 ;
      LAYER Metal4 ;
        RECT 152.17 12 152.83 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 176.33 12 176.99 12.66 ;
      LAYER Metal6 ;
        RECT 176.33 12 176.99 12.66 ;
      LAYER Metal3 ;
        RECT 176.33 12 176.99 12.66 ;
      LAYER Metal4 ;
        RECT 176.33 12 176.99 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 194.73 12 195.39 12.66 ;
      LAYER Metal6 ;
        RECT 194.73 12 195.39 12.66 ;
      LAYER Metal3 ;
        RECT 194.73 12 195.39 12.66 ;
      LAYER Metal4 ;
        RECT 194.73 12 195.39 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.89 12 219.55 12.66 ;
      LAYER Metal6 ;
        RECT 218.89 12 219.55 12.66 ;
      LAYER Metal3 ;
        RECT 218.89 12 219.55 12.66 ;
      LAYER Metal4 ;
        RECT 218.89 12 219.55 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 27.37 12 28.03 12.66 ;
      LAYER Metal6 ;
        RECT 27.37 12 28.03 12.66 ;
      LAYER Metal3 ;
        RECT 27.37 12 28.03 12.66 ;
      LAYER Metal4 ;
        RECT 27.37 12 28.03 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 240.17 12 240.83 12.66 ;
      LAYER Metal6 ;
        RECT 240.17 12 240.83 12.66 ;
      LAYER Metal3 ;
        RECT 240.17 12 240.83 12.66 ;
      LAYER Metal4 ;
        RECT 240.17 12 240.83 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 258.57 12 259.23 12.66 ;
      LAYER Metal6 ;
        RECT 258.57 12 259.23 12.66 ;
      LAYER Metal3 ;
        RECT 258.57 12 259.23 12.66 ;
      LAYER Metal4 ;
        RECT 258.57 12 259.23 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 282.73 12 283.39 12.66 ;
      LAYER Metal6 ;
        RECT 282.73 12 283.39 12.66 ;
      LAYER Metal3 ;
        RECT 282.73 12 283.39 12.66 ;
      LAYER Metal4 ;
        RECT 282.73 12 283.39 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 301.13 12 301.79 12.66 ;
      LAYER Metal6 ;
        RECT 301.13 12 301.79 12.66 ;
      LAYER Metal3 ;
        RECT 301.13 12 301.79 12.66 ;
      LAYER Metal4 ;
        RECT 301.13 12 301.79 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 325.29 12 325.95 12.66 ;
      LAYER Metal6 ;
        RECT 325.29 12 325.95 12.66 ;
      LAYER Metal3 ;
        RECT 325.29 12 325.95 12.66 ;
      LAYER Metal4 ;
        RECT 325.29 12 325.95 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 343.69 12 344.35 12.66 ;
      LAYER Metal6 ;
        RECT 343.69 12 344.35 12.66 ;
      LAYER Metal3 ;
        RECT 343.69 12 344.35 12.66 ;
      LAYER Metal4 ;
        RECT 343.69 12 344.35 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 404.935 12 405.595 12.66 ;
      LAYER Metal6 ;
        RECT 404.935 12 405.595 12.66 ;
      LAYER Metal3 ;
        RECT 404.935 12 405.595 12.66 ;
      LAYER Metal4 ;
        RECT 404.935 12 405.595 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 423.335 12 423.995 12.66 ;
      LAYER Metal6 ;
        RECT 423.335 12 423.995 12.66 ;
      LAYER Metal3 ;
        RECT 423.335 12 423.995 12.66 ;
      LAYER Metal4 ;
        RECT 423.335 12 423.995 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 447.495 12 448.155 12.66 ;
      LAYER Metal6 ;
        RECT 447.495 12 448.155 12.66 ;
      LAYER Metal3 ;
        RECT 447.495 12 448.155 12.66 ;
      LAYER Metal4 ;
        RECT 447.495 12 448.155 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 465.895 12 466.555 12.66 ;
      LAYER Metal6 ;
        RECT 465.895 12 466.555 12.66 ;
      LAYER Metal3 ;
        RECT 465.895 12 466.555 12.66 ;
      LAYER Metal4 ;
        RECT 465.895 12 466.555 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 45.77 12 46.43 12.66 ;
      LAYER Metal6 ;
        RECT 45.77 12 46.43 12.66 ;
      LAYER Metal3 ;
        RECT 45.77 12 46.43 12.66 ;
      LAYER Metal4 ;
        RECT 45.77 12 46.43 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 490.055 12 490.715 12.66 ;
      LAYER Metal6 ;
        RECT 490.055 12 490.715 12.66 ;
      LAYER Metal3 ;
        RECT 490.055 12 490.715 12.66 ;
      LAYER Metal4 ;
        RECT 490.055 12 490.715 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 508.455 12 509.115 12.66 ;
      LAYER Metal6 ;
        RECT 508.455 12 509.115 12.66 ;
      LAYER Metal3 ;
        RECT 508.455 12 509.115 12.66 ;
      LAYER Metal4 ;
        RECT 508.455 12 509.115 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 532.615 12 533.275 12.66 ;
      LAYER Metal6 ;
        RECT 532.615 12 533.275 12.66 ;
      LAYER Metal3 ;
        RECT 532.615 12 533.275 12.66 ;
      LAYER Metal4 ;
        RECT 532.615 12 533.275 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 551.015 12 551.675 12.66 ;
      LAYER Metal6 ;
        RECT 551.015 12 551.675 12.66 ;
      LAYER Metal3 ;
        RECT 551.015 12 551.675 12.66 ;
      LAYER Metal4 ;
        RECT 551.015 12 551.675 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 575.175 12 575.835 12.66 ;
      LAYER Metal6 ;
        RECT 575.175 12 575.835 12.66 ;
      LAYER Metal3 ;
        RECT 575.175 12 575.835 12.66 ;
      LAYER Metal4 ;
        RECT 575.175 12 575.835 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 593.575 12 594.235 12.66 ;
      LAYER Metal6 ;
        RECT 593.575 12 594.235 12.66 ;
      LAYER Metal3 ;
        RECT 593.575 12 594.235 12.66 ;
      LAYER Metal4 ;
        RECT 593.575 12 594.235 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 617.735 12 618.395 12.66 ;
      LAYER Metal6 ;
        RECT 617.735 12 618.395 12.66 ;
      LAYER Metal3 ;
        RECT 617.735 12 618.395 12.66 ;
      LAYER Metal4 ;
        RECT 617.735 12 618.395 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 636.135 12 636.795 12.66 ;
      LAYER Metal6 ;
        RECT 636.135 12 636.795 12.66 ;
      LAYER Metal3 ;
        RECT 636.135 12 636.795 12.66 ;
      LAYER Metal4 ;
        RECT 636.135 12 636.795 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 660.295 12 660.955 12.66 ;
      LAYER Metal6 ;
        RECT 660.295 12 660.955 12.66 ;
      LAYER Metal3 ;
        RECT 660.295 12 660.955 12.66 ;
      LAYER Metal4 ;
        RECT 660.295 12 660.955 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 678.695 12 679.355 12.66 ;
      LAYER Metal6 ;
        RECT 678.695 12 679.355 12.66 ;
      LAYER Metal3 ;
        RECT 678.695 12 679.355 12.66 ;
      LAYER Metal4 ;
        RECT 678.695 12 679.355 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.93 12 70.59 12.66 ;
      LAYER Metal6 ;
        RECT 69.93 12 70.59 12.66 ;
      LAYER Metal3 ;
        RECT 69.93 12 70.59 12.66 ;
      LAYER Metal4 ;
        RECT 69.93 12 70.59 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 702.855 12 703.515 12.66 ;
      LAYER Metal6 ;
        RECT 702.855 12 703.515 12.66 ;
      LAYER Metal3 ;
        RECT 702.855 12 703.515 12.66 ;
      LAYER Metal4 ;
        RECT 702.855 12 703.515 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 721.255 12 721.915 12.66 ;
      LAYER Metal6 ;
        RECT 721.255 12 721.915 12.66 ;
      LAYER Metal3 ;
        RECT 721.255 12 721.915 12.66 ;
      LAYER Metal4 ;
        RECT 721.255 12 721.915 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 88.33 12 88.99 12.66 ;
      LAYER Metal6 ;
        RECT 88.33 12 88.99 12.66 ;
      LAYER Metal3 ;
        RECT 88.33 12 88.99 12.66 ;
      LAYER Metal4 ;
        RECT 88.33 12 88.99 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 112.49 12 113.15 12.66 ;
      LAYER Metal6 ;
        RECT 112.49 12 113.15 12.66 ;
      LAYER Metal3 ;
        RECT 112.49 12 113.15 12.66 ;
      LAYER Metal4 ;
        RECT 112.49 12 113.15 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 130.89 12 131.55 12.66 ;
      LAYER Metal6 ;
        RECT 130.89 12 131.55 12.66 ;
      LAYER Metal3 ;
        RECT 130.89 12 131.55 12.66 ;
      LAYER Metal4 ;
        RECT 130.89 12 131.55 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 155.05 12 155.71 12.66 ;
      LAYER Metal6 ;
        RECT 155.05 12 155.71 12.66 ;
      LAYER Metal3 ;
        RECT 155.05 12 155.71 12.66 ;
      LAYER Metal4 ;
        RECT 155.05 12 155.71 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 173.45 12 174.11 12.66 ;
      LAYER Metal6 ;
        RECT 173.45 12 174.11 12.66 ;
      LAYER Metal3 ;
        RECT 173.45 12 174.11 12.66 ;
      LAYER Metal4 ;
        RECT 173.45 12 174.11 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 197.61 12 198.27 12.66 ;
      LAYER Metal6 ;
        RECT 197.61 12 198.27 12.66 ;
      LAYER Metal3 ;
        RECT 197.61 12 198.27 12.66 ;
      LAYER Metal4 ;
        RECT 197.61 12 198.27 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 216.01 12 216.67 12.66 ;
      LAYER Metal6 ;
        RECT 216.01 12 216.67 12.66 ;
      LAYER Metal3 ;
        RECT 216.01 12 216.67 12.66 ;
      LAYER Metal4 ;
        RECT 216.01 12 216.67 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.425 12 385.085 12.66 ;
      LAYER Metal6 ;
        RECT 384.425 12 385.085 12.66 ;
      LAYER Metal3 ;
        RECT 384.425 12 385.085 12.66 ;
      LAYER Metal4 ;
        RECT 384.425 12 385.085 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 364.2 12 364.86 12.66 ;
      LAYER Metal6 ;
        RECT 364.2 12 364.86 12.66 ;
      LAYER Metal3 ;
        RECT 364.2 12 364.86 12.66 ;
      LAYER Metal4 ;
        RECT 364.2 12 364.86 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 302.3 772.885 307.3 ;
        RECT 0 0 772.885 5 ;
      LAYER Metal2 ;
        RECT 0 0 5 307.3 ;
        RECT 767.885 0 772.885 307.3 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 296.7 767.285 301.7 ;
        RECT 5.6 5.6 767.285 10.6 ;
      LAYER Metal2 ;
        RECT 5.6 5.6 10.6 301.7 ;
        RECT 762.285 5.6 767.285 301.7 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 760.88 295.255 ;
    LAYER Metal2 ;
      RECT 12 12 760.88 295.255 ;
    LAYER Metal3 ;
      RECT 12 12 760.88 295.255 ;
    LAYER Metal4 ;
      RECT 12 12 760.88 295.255 ;
    LAYER Metal5 ;
      RECT 12 12 760.88 295.255 ;
    LAYER Metal6 ;
      RECT 12 12 760.88 295.255 ;
  END
END MEM2_1024X32

END LIBRARY
