VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MEM2_128X32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2_128X32 0 0 ;
  SIZE 423.015 BY 145.035 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 102.42 12.66 103.08 ;
      LAYER Metal6 ;
        RECT 12 102.42 12.66 103.08 ;
      LAYER Metal3 ;
        RECT 12 102.42 12.66 103.08 ;
      LAYER Metal4 ;
        RECT 12 102.42 12.66 103.08 ;
    END
  END A1[0]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 96.3 12.66 96.96 ;
      LAYER Metal6 ;
        RECT 12 96.3 12.66 96.96 ;
      LAYER Metal3 ;
        RECT 12 96.3 12.66 96.96 ;
      LAYER Metal4 ;
        RECT 12 96.3 12.66 96.96 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 87.08 12.66 87.74 ;
      LAYER Metal6 ;
        RECT 12 87.08 12.66 87.74 ;
      LAYER Metal3 ;
        RECT 12 87.08 12.66 87.74 ;
      LAYER Metal4 ;
        RECT 12 87.08 12.66 87.74 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 84.06 12.66 84.72 ;
      LAYER Metal6 ;
        RECT 12 84.06 12.66 84.72 ;
      LAYER Metal3 ;
        RECT 12 84.06 12.66 84.72 ;
      LAYER Metal4 ;
        RECT 12 84.06 12.66 84.72 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 80.96 12.66 81.62 ;
      LAYER Metal6 ;
        RECT 12 80.96 12.66 81.62 ;
      LAYER Metal3 ;
        RECT 12 80.96 12.66 81.62 ;
      LAYER Metal4 ;
        RECT 12 80.96 12.66 81.62 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 74.84 12.66 75.5 ;
      LAYER Metal6 ;
        RECT 12 74.84 12.66 75.5 ;
      LAYER Metal3 ;
        RECT 12 74.84 12.66 75.5 ;
      LAYER Metal4 ;
        RECT 12 74.84 12.66 75.5 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 71.82 12.66 72.48 ;
      LAYER Metal6 ;
        RECT 12 71.82 12.66 72.48 ;
      LAYER Metal3 ;
        RECT 12 71.82 12.66 72.48 ;
      LAYER Metal4 ;
        RECT 12 71.82 12.66 72.48 ;
    END
  END A1[6]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 36.4 12.66 37.06 ;
      LAYER Metal6 ;
        RECT 12 36.4 12.66 37.06 ;
      LAYER Metal3 ;
        RECT 12 36.4 12.66 37.06 ;
      LAYER Metal4 ;
        RECT 12 36.4 12.66 37.06 ;
    END
  END A2[0]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 42.52 12.66 43.18 ;
      LAYER Metal6 ;
        RECT 12 42.52 12.66 43.18 ;
      LAYER Metal3 ;
        RECT 12 42.52 12.66 43.18 ;
      LAYER Metal4 ;
        RECT 12 42.52 12.66 43.18 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 51.74 12.66 52.4 ;
      LAYER Metal6 ;
        RECT 12 51.74 12.66 52.4 ;
      LAYER Metal3 ;
        RECT 12 51.74 12.66 52.4 ;
      LAYER Metal4 ;
        RECT 12 51.74 12.66 52.4 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 54.76 12.66 55.42 ;
      LAYER Metal6 ;
        RECT 12 54.76 12.66 55.42 ;
      LAYER Metal3 ;
        RECT 12 54.76 12.66 55.42 ;
      LAYER Metal4 ;
        RECT 12 54.76 12.66 55.42 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 57.86 12.66 58.52 ;
      LAYER Metal6 ;
        RECT 12 57.86 12.66 58.52 ;
      LAYER Metal3 ;
        RECT 12 57.86 12.66 58.52 ;
      LAYER Metal4 ;
        RECT 12 57.86 12.66 58.52 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 63.98 12.66 64.64 ;
      LAYER Metal6 ;
        RECT 12 63.98 12.66 64.64 ;
      LAYER Metal3 ;
        RECT 12 63.98 12.66 64.64 ;
      LAYER Metal4 ;
        RECT 12 63.98 12.66 64.64 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 67 12.66 67.66 ;
      LAYER Metal6 ;
        RECT 12 67 12.66 67.66 ;
      LAYER Metal3 ;
        RECT 12 67 12.66 67.66 ;
      LAYER Metal4 ;
        RECT 12 67 12.66 67.66 ;
    END
  END A2[6]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 210.28 12 210.94 12.66 ;
      LAYER Metal6 ;
        RECT 210.28 12 210.94 12.66 ;
      LAYER Metal3 ;
        RECT 210.28 12 210.94 12.66 ;
      LAYER Metal4 ;
        RECT 210.28 12 210.94 12.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal6 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal3 ;
        RECT 196.36 12 197.02 12.66 ;
      LAYER Metal4 ;
        RECT 196.36 12 197.02 12.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 218.905 12 219.565 12.66 ;
      LAYER Metal6 ;
        RECT 218.905 12 219.565 12.66 ;
      LAYER Metal3 ;
        RECT 218.905 12 219.565 12.66 ;
      LAYER Metal4 ;
        RECT 218.905 12 219.565 12.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal6 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal3 ;
        RECT 187.735 12 188.395 12.66 ;
      LAYER Metal4 ;
        RECT 187.735 12 188.395 12.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal6 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal3 ;
        RECT 15.86 12 16.52 12.66 ;
      LAYER Metal4 ;
        RECT 15.86 12 16.52 12.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal6 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal3 ;
        RECT 122.26 12 122.92 12.66 ;
      LAYER Metal4 ;
        RECT 122.26 12 122.92 12.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal6 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal3 ;
        RECT 142.4 12 143.06 12.66 ;
      LAYER Metal4 ;
        RECT 142.4 12 143.06 12.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal6 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal3 ;
        RECT 143.54 12 144.2 12.66 ;
      LAYER Metal4 ;
        RECT 143.54 12 144.2 12.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal6 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal3 ;
        RECT 163.68 12 164.34 12.66 ;
      LAYER Metal4 ;
        RECT 163.68 12 164.34 12.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal6 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal3 ;
        RECT 164.82 12 165.48 12.66 ;
      LAYER Metal4 ;
        RECT 164.82 12 165.48 12.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal6 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal3 ;
        RECT 184.96 12 185.62 12.66 ;
      LAYER Metal4 ;
        RECT 184.96 12 185.62 12.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 221.68 12 222.34 12.66 ;
      LAYER Metal6 ;
        RECT 221.68 12 222.34 12.66 ;
      LAYER Metal3 ;
        RECT 221.68 12 222.34 12.66 ;
      LAYER Metal4 ;
        RECT 221.68 12 222.34 12.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 241.82 12 242.48 12.66 ;
      LAYER Metal6 ;
        RECT 241.82 12 242.48 12.66 ;
      LAYER Metal3 ;
        RECT 241.82 12 242.48 12.66 ;
      LAYER Metal4 ;
        RECT 241.82 12 242.48 12.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 242.96 12 243.62 12.66 ;
      LAYER Metal6 ;
        RECT 242.96 12 243.62 12.66 ;
      LAYER Metal3 ;
        RECT 242.96 12 243.62 12.66 ;
      LAYER Metal4 ;
        RECT 242.96 12 243.62 12.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 263.1 12 263.76 12.66 ;
      LAYER Metal6 ;
        RECT 263.1 12 263.76 12.66 ;
      LAYER Metal3 ;
        RECT 263.1 12 263.76 12.66 ;
      LAYER Metal4 ;
        RECT 263.1 12 263.76 12.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal6 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal3 ;
        RECT 36 12 36.66 12.66 ;
      LAYER Metal4 ;
        RECT 36 12 36.66 12.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 264.24 12 264.9 12.66 ;
      LAYER Metal6 ;
        RECT 264.24 12 264.9 12.66 ;
      LAYER Metal3 ;
        RECT 264.24 12 264.9 12.66 ;
      LAYER Metal4 ;
        RECT 264.24 12 264.9 12.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 284.38 12 285.04 12.66 ;
      LAYER Metal6 ;
        RECT 284.38 12 285.04 12.66 ;
      LAYER Metal3 ;
        RECT 284.38 12 285.04 12.66 ;
      LAYER Metal4 ;
        RECT 284.38 12 285.04 12.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 285.52 12 286.18 12.66 ;
      LAYER Metal6 ;
        RECT 285.52 12 286.18 12.66 ;
      LAYER Metal3 ;
        RECT 285.52 12 286.18 12.66 ;
      LAYER Metal4 ;
        RECT 285.52 12 286.18 12.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 305.66 12 306.32 12.66 ;
      LAYER Metal6 ;
        RECT 305.66 12 306.32 12.66 ;
      LAYER Metal3 ;
        RECT 305.66 12 306.32 12.66 ;
      LAYER Metal4 ;
        RECT 305.66 12 306.32 12.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.8 12 307.46 12.66 ;
      LAYER Metal6 ;
        RECT 306.8 12 307.46 12.66 ;
      LAYER Metal3 ;
        RECT 306.8 12 307.46 12.66 ;
      LAYER Metal4 ;
        RECT 306.8 12 307.46 12.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 326.94 12 327.6 12.66 ;
      LAYER Metal6 ;
        RECT 326.94 12 327.6 12.66 ;
      LAYER Metal3 ;
        RECT 326.94 12 327.6 12.66 ;
      LAYER Metal4 ;
        RECT 326.94 12 327.6 12.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 328.08 12 328.74 12.66 ;
      LAYER Metal6 ;
        RECT 328.08 12 328.74 12.66 ;
      LAYER Metal3 ;
        RECT 328.08 12 328.74 12.66 ;
      LAYER Metal4 ;
        RECT 328.08 12 328.74 12.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 348.22 12 348.88 12.66 ;
      LAYER Metal6 ;
        RECT 348.22 12 348.88 12.66 ;
      LAYER Metal3 ;
        RECT 348.22 12 348.88 12.66 ;
      LAYER Metal4 ;
        RECT 348.22 12 348.88 12.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 349.36 12 350.02 12.66 ;
      LAYER Metal6 ;
        RECT 349.36 12 350.02 12.66 ;
      LAYER Metal3 ;
        RECT 349.36 12 350.02 12.66 ;
      LAYER Metal4 ;
        RECT 349.36 12 350.02 12.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 369.5 12 370.16 12.66 ;
      LAYER Metal6 ;
        RECT 369.5 12 370.16 12.66 ;
      LAYER Metal3 ;
        RECT 369.5 12 370.16 12.66 ;
      LAYER Metal4 ;
        RECT 369.5 12 370.16 12.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal6 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal3 ;
        RECT 37.14 12 37.8 12.66 ;
      LAYER Metal4 ;
        RECT 37.14 12 37.8 12.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 370.64 12 371.3 12.66 ;
      LAYER Metal6 ;
        RECT 370.64 12 371.3 12.66 ;
      LAYER Metal3 ;
        RECT 370.64 12 371.3 12.66 ;
      LAYER Metal4 ;
        RECT 370.64 12 371.3 12.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 390.78 12 391.44 12.66 ;
      LAYER Metal6 ;
        RECT 390.78 12 391.44 12.66 ;
      LAYER Metal3 ;
        RECT 390.78 12 391.44 12.66 ;
      LAYER Metal4 ;
        RECT 390.78 12 391.44 12.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal6 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal3 ;
        RECT 57.28 12 57.94 12.66 ;
      LAYER Metal4 ;
        RECT 57.28 12 57.94 12.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal6 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal3 ;
        RECT 58.42 12 59.08 12.66 ;
      LAYER Metal4 ;
        RECT 58.42 12 59.08 12.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal6 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal3 ;
        RECT 78.56 12 79.22 12.66 ;
      LAYER Metal4 ;
        RECT 78.56 12 79.22 12.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal6 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal3 ;
        RECT 79.7 12 80.36 12.66 ;
      LAYER Metal4 ;
        RECT 79.7 12 80.36 12.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal6 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal3 ;
        RECT 99.84 12 100.5 12.66 ;
      LAYER Metal4 ;
        RECT 99.84 12 100.5 12.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal6 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal3 ;
        RECT 100.98 12 101.64 12.66 ;
      LAYER Metal4 ;
        RECT 100.98 12 101.64 12.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal6 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal3 ;
        RECT 121.12 12 121.78 12.66 ;
      LAYER Metal4 ;
        RECT 121.12 12 121.78 12.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal6 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal3 ;
        RECT 25.36 12 26.02 12.66 ;
      LAYER Metal4 ;
        RECT 25.36 12 26.02 12.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal6 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal3 ;
        RECT 131.76 12 132.42 12.66 ;
      LAYER Metal4 ;
        RECT 131.76 12 132.42 12.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal6 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal3 ;
        RECT 132.9 12 133.56 12.66 ;
      LAYER Metal4 ;
        RECT 132.9 12 133.56 12.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal6 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal3 ;
        RECT 153.04 12 153.7 12.66 ;
      LAYER Metal4 ;
        RECT 153.04 12 153.7 12.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal6 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal3 ;
        RECT 154.18 12 154.84 12.66 ;
      LAYER Metal4 ;
        RECT 154.18 12 154.84 12.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal6 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal3 ;
        RECT 174.32 12 174.98 12.66 ;
      LAYER Metal4 ;
        RECT 174.32 12 174.98 12.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal6 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal3 ;
        RECT 175.46 12 176.12 12.66 ;
      LAYER Metal4 ;
        RECT 175.46 12 176.12 12.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 231.18 12 231.84 12.66 ;
      LAYER Metal6 ;
        RECT 231.18 12 231.84 12.66 ;
      LAYER Metal3 ;
        RECT 231.18 12 231.84 12.66 ;
      LAYER Metal4 ;
        RECT 231.18 12 231.84 12.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 232.32 12 232.98 12.66 ;
      LAYER Metal6 ;
        RECT 232.32 12 232.98 12.66 ;
      LAYER Metal3 ;
        RECT 232.32 12 232.98 12.66 ;
      LAYER Metal4 ;
        RECT 232.32 12 232.98 12.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 252.46 12 253.12 12.66 ;
      LAYER Metal6 ;
        RECT 252.46 12 253.12 12.66 ;
      LAYER Metal3 ;
        RECT 252.46 12 253.12 12.66 ;
      LAYER Metal4 ;
        RECT 252.46 12 253.12 12.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 253.6 12 254.26 12.66 ;
      LAYER Metal6 ;
        RECT 253.6 12 254.26 12.66 ;
      LAYER Metal3 ;
        RECT 253.6 12 254.26 12.66 ;
      LAYER Metal4 ;
        RECT 253.6 12 254.26 12.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal6 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal3 ;
        RECT 26.5 12 27.16 12.66 ;
      LAYER Metal4 ;
        RECT 26.5 12 27.16 12.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 273.74 12 274.4 12.66 ;
      LAYER Metal6 ;
        RECT 273.74 12 274.4 12.66 ;
      LAYER Metal3 ;
        RECT 273.74 12 274.4 12.66 ;
      LAYER Metal4 ;
        RECT 273.74 12 274.4 12.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 274.88 12 275.54 12.66 ;
      LAYER Metal6 ;
        RECT 274.88 12 275.54 12.66 ;
      LAYER Metal3 ;
        RECT 274.88 12 275.54 12.66 ;
      LAYER Metal4 ;
        RECT 274.88 12 275.54 12.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 295.02 12 295.68 12.66 ;
      LAYER Metal6 ;
        RECT 295.02 12 295.68 12.66 ;
      LAYER Metal3 ;
        RECT 295.02 12 295.68 12.66 ;
      LAYER Metal4 ;
        RECT 295.02 12 295.68 12.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 296.16 12 296.82 12.66 ;
      LAYER Metal6 ;
        RECT 296.16 12 296.82 12.66 ;
      LAYER Metal3 ;
        RECT 296.16 12 296.82 12.66 ;
      LAYER Metal4 ;
        RECT 296.16 12 296.82 12.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 316.3 12 316.96 12.66 ;
      LAYER Metal6 ;
        RECT 316.3 12 316.96 12.66 ;
      LAYER Metal3 ;
        RECT 316.3 12 316.96 12.66 ;
      LAYER Metal4 ;
        RECT 316.3 12 316.96 12.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 317.44 12 318.1 12.66 ;
      LAYER Metal6 ;
        RECT 317.44 12 318.1 12.66 ;
      LAYER Metal3 ;
        RECT 317.44 12 318.1 12.66 ;
      LAYER Metal4 ;
        RECT 317.44 12 318.1 12.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 337.58 12 338.24 12.66 ;
      LAYER Metal6 ;
        RECT 337.58 12 338.24 12.66 ;
      LAYER Metal3 ;
        RECT 337.58 12 338.24 12.66 ;
      LAYER Metal4 ;
        RECT 337.58 12 338.24 12.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 338.72 12 339.38 12.66 ;
      LAYER Metal6 ;
        RECT 338.72 12 339.38 12.66 ;
      LAYER Metal3 ;
        RECT 338.72 12 339.38 12.66 ;
      LAYER Metal4 ;
        RECT 338.72 12 339.38 12.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 358.86 12 359.52 12.66 ;
      LAYER Metal6 ;
        RECT 358.86 12 359.52 12.66 ;
      LAYER Metal3 ;
        RECT 358.86 12 359.52 12.66 ;
      LAYER Metal4 ;
        RECT 358.86 12 359.52 12.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 360 12 360.66 12.66 ;
      LAYER Metal6 ;
        RECT 360 12 360.66 12.66 ;
      LAYER Metal3 ;
        RECT 360 12 360.66 12.66 ;
      LAYER Metal4 ;
        RECT 360 12 360.66 12.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal6 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal3 ;
        RECT 46.64 12 47.3 12.66 ;
      LAYER Metal4 ;
        RECT 46.64 12 47.3 12.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 380.14 12 380.8 12.66 ;
      LAYER Metal6 ;
        RECT 380.14 12 380.8 12.66 ;
      LAYER Metal3 ;
        RECT 380.14 12 380.8 12.66 ;
      LAYER Metal4 ;
        RECT 380.14 12 380.8 12.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 381.28 12 381.94 12.66 ;
      LAYER Metal6 ;
        RECT 381.28 12 381.94 12.66 ;
      LAYER Metal3 ;
        RECT 381.28 12 381.94 12.66 ;
      LAYER Metal4 ;
        RECT 381.28 12 381.94 12.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal6 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal3 ;
        RECT 47.78 12 48.44 12.66 ;
      LAYER Metal4 ;
        RECT 47.78 12 48.44 12.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal6 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal3 ;
        RECT 67.92 12 68.58 12.66 ;
      LAYER Metal4 ;
        RECT 67.92 12 68.58 12.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal6 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal3 ;
        RECT 69.06 12 69.72 12.66 ;
      LAYER Metal4 ;
        RECT 69.06 12 69.72 12.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal6 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal3 ;
        RECT 89.2 12 89.86 12.66 ;
      LAYER Metal4 ;
        RECT 89.2 12 89.86 12.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal6 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal3 ;
        RECT 90.34 12 91 12.66 ;
      LAYER Metal4 ;
        RECT 90.34 12 91 12.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal6 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal3 ;
        RECT 110.48 12 111.14 12.66 ;
      LAYER Metal4 ;
        RECT 110.48 12 111.14 12.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal6 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal3 ;
        RECT 111.62 12 112.28 12.66 ;
      LAYER Metal4 ;
        RECT 111.62 12 112.28 12.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal6 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal3 ;
        RECT 18.28 12 18.94 12.66 ;
      LAYER Metal4 ;
        RECT 18.28 12 18.94 12.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal6 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal3 ;
        RECT 125.56 12 126.22 12.66 ;
      LAYER Metal4 ;
        RECT 125.56 12 126.22 12.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal6 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal3 ;
        RECT 139.1 12 139.76 12.66 ;
      LAYER Metal4 ;
        RECT 139.1 12 139.76 12.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal6 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal3 ;
        RECT 146.84 12 147.5 12.66 ;
      LAYER Metal4 ;
        RECT 146.84 12 147.5 12.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal6 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal3 ;
        RECT 160.38 12 161.04 12.66 ;
      LAYER Metal4 ;
        RECT 160.38 12 161.04 12.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal6 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal3 ;
        RECT 168.12 12 168.78 12.66 ;
      LAYER Metal4 ;
        RECT 168.12 12 168.78 12.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal6 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal3 ;
        RECT 181.66 12 182.32 12.66 ;
      LAYER Metal4 ;
        RECT 181.66 12 182.32 12.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 224.98 12 225.64 12.66 ;
      LAYER Metal6 ;
        RECT 224.98 12 225.64 12.66 ;
      LAYER Metal3 ;
        RECT 224.98 12 225.64 12.66 ;
      LAYER Metal4 ;
        RECT 224.98 12 225.64 12.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 238.52 12 239.18 12.66 ;
      LAYER Metal6 ;
        RECT 238.52 12 239.18 12.66 ;
      LAYER Metal3 ;
        RECT 238.52 12 239.18 12.66 ;
      LAYER Metal4 ;
        RECT 238.52 12 239.18 12.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 246.26 12 246.92 12.66 ;
      LAYER Metal6 ;
        RECT 246.26 12 246.92 12.66 ;
      LAYER Metal3 ;
        RECT 246.26 12 246.92 12.66 ;
      LAYER Metal4 ;
        RECT 246.26 12 246.92 12.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 259.8 12 260.46 12.66 ;
      LAYER Metal6 ;
        RECT 259.8 12 260.46 12.66 ;
      LAYER Metal3 ;
        RECT 259.8 12 260.46 12.66 ;
      LAYER Metal4 ;
        RECT 259.8 12 260.46 12.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal6 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal3 ;
        RECT 32.7 12 33.36 12.66 ;
      LAYER Metal4 ;
        RECT 32.7 12 33.36 12.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 267.54 12 268.2 12.66 ;
      LAYER Metal6 ;
        RECT 267.54 12 268.2 12.66 ;
      LAYER Metal3 ;
        RECT 267.54 12 268.2 12.66 ;
      LAYER Metal4 ;
        RECT 267.54 12 268.2 12.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 281.08 12 281.74 12.66 ;
      LAYER Metal6 ;
        RECT 281.08 12 281.74 12.66 ;
      LAYER Metal3 ;
        RECT 281.08 12 281.74 12.66 ;
      LAYER Metal4 ;
        RECT 281.08 12 281.74 12.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 288.82 12 289.48 12.66 ;
      LAYER Metal6 ;
        RECT 288.82 12 289.48 12.66 ;
      LAYER Metal3 ;
        RECT 288.82 12 289.48 12.66 ;
      LAYER Metal4 ;
        RECT 288.82 12 289.48 12.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 302.36 12 303.02 12.66 ;
      LAYER Metal6 ;
        RECT 302.36 12 303.02 12.66 ;
      LAYER Metal3 ;
        RECT 302.36 12 303.02 12.66 ;
      LAYER Metal4 ;
        RECT 302.36 12 303.02 12.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 310.1 12 310.76 12.66 ;
      LAYER Metal6 ;
        RECT 310.1 12 310.76 12.66 ;
      LAYER Metal3 ;
        RECT 310.1 12 310.76 12.66 ;
      LAYER Metal4 ;
        RECT 310.1 12 310.76 12.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 323.64 12 324.3 12.66 ;
      LAYER Metal6 ;
        RECT 323.64 12 324.3 12.66 ;
      LAYER Metal3 ;
        RECT 323.64 12 324.3 12.66 ;
      LAYER Metal4 ;
        RECT 323.64 12 324.3 12.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 331.38 12 332.04 12.66 ;
      LAYER Metal6 ;
        RECT 331.38 12 332.04 12.66 ;
      LAYER Metal3 ;
        RECT 331.38 12 332.04 12.66 ;
      LAYER Metal4 ;
        RECT 331.38 12 332.04 12.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 344.92 12 345.58 12.66 ;
      LAYER Metal6 ;
        RECT 344.92 12 345.58 12.66 ;
      LAYER Metal3 ;
        RECT 344.92 12 345.58 12.66 ;
      LAYER Metal4 ;
        RECT 344.92 12 345.58 12.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 352.66 12 353.32 12.66 ;
      LAYER Metal6 ;
        RECT 352.66 12 353.32 12.66 ;
      LAYER Metal3 ;
        RECT 352.66 12 353.32 12.66 ;
      LAYER Metal4 ;
        RECT 352.66 12 353.32 12.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 366.2 12 366.86 12.66 ;
      LAYER Metal6 ;
        RECT 366.2 12 366.86 12.66 ;
      LAYER Metal3 ;
        RECT 366.2 12 366.86 12.66 ;
      LAYER Metal4 ;
        RECT 366.2 12 366.86 12.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal6 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal3 ;
        RECT 40.44 12 41.1 12.66 ;
      LAYER Metal4 ;
        RECT 40.44 12 41.1 12.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 373.94 12 374.6 12.66 ;
      LAYER Metal6 ;
        RECT 373.94 12 374.6 12.66 ;
      LAYER Metal3 ;
        RECT 373.94 12 374.6 12.66 ;
      LAYER Metal4 ;
        RECT 373.94 12 374.6 12.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 388.36 12 389.02 12.66 ;
      LAYER Metal6 ;
        RECT 388.36 12 389.02 12.66 ;
      LAYER Metal3 ;
        RECT 388.36 12 389.02 12.66 ;
      LAYER Metal4 ;
        RECT 388.36 12 389.02 12.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal6 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal3 ;
        RECT 53.98 12 54.64 12.66 ;
      LAYER Metal4 ;
        RECT 53.98 12 54.64 12.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal6 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal3 ;
        RECT 61.72 12 62.38 12.66 ;
      LAYER Metal4 ;
        RECT 61.72 12 62.38 12.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal6 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal3 ;
        RECT 75.26 12 75.92 12.66 ;
      LAYER Metal4 ;
        RECT 75.26 12 75.92 12.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal6 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal3 ;
        RECT 83 12 83.66 12.66 ;
      LAYER Metal4 ;
        RECT 83 12 83.66 12.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal6 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal3 ;
        RECT 96.54 12 97.2 12.66 ;
      LAYER Metal4 ;
        RECT 96.54 12 97.2 12.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal6 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal3 ;
        RECT 104.28 12 104.94 12.66 ;
      LAYER Metal4 ;
        RECT 104.28 12 104.94 12.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal6 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal3 ;
        RECT 117.82 12 118.48 12.66 ;
      LAYER Metal4 ;
        RECT 117.82 12 118.48 12.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal6 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal3 ;
        RECT 22.06 12 22.72 12.66 ;
      LAYER Metal4 ;
        RECT 22.06 12 22.72 12.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal6 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal3 ;
        RECT 128.46 12 129.12 12.66 ;
      LAYER Metal4 ;
        RECT 128.46 12 129.12 12.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal6 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal3 ;
        RECT 136.2 12 136.86 12.66 ;
      LAYER Metal4 ;
        RECT 136.2 12 136.86 12.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal6 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal3 ;
        RECT 149.74 12 150.4 12.66 ;
      LAYER Metal4 ;
        RECT 149.74 12 150.4 12.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal6 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal3 ;
        RECT 157.48 12 158.14 12.66 ;
      LAYER Metal4 ;
        RECT 157.48 12 158.14 12.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal6 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal3 ;
        RECT 171.02 12 171.68 12.66 ;
      LAYER Metal4 ;
        RECT 171.02 12 171.68 12.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal6 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal3 ;
        RECT 178.76 12 179.42 12.66 ;
      LAYER Metal4 ;
        RECT 178.76 12 179.42 12.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 227.88 12 228.54 12.66 ;
      LAYER Metal6 ;
        RECT 227.88 12 228.54 12.66 ;
      LAYER Metal3 ;
        RECT 227.88 12 228.54 12.66 ;
      LAYER Metal4 ;
        RECT 227.88 12 228.54 12.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 235.62 12 236.28 12.66 ;
      LAYER Metal6 ;
        RECT 235.62 12 236.28 12.66 ;
      LAYER Metal3 ;
        RECT 235.62 12 236.28 12.66 ;
      LAYER Metal4 ;
        RECT 235.62 12 236.28 12.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 249.16 12 249.82 12.66 ;
      LAYER Metal6 ;
        RECT 249.16 12 249.82 12.66 ;
      LAYER Metal3 ;
        RECT 249.16 12 249.82 12.66 ;
      LAYER Metal4 ;
        RECT 249.16 12 249.82 12.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 256.9 12 257.56 12.66 ;
      LAYER Metal6 ;
        RECT 256.9 12 257.56 12.66 ;
      LAYER Metal3 ;
        RECT 256.9 12 257.56 12.66 ;
      LAYER Metal4 ;
        RECT 256.9 12 257.56 12.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal6 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal3 ;
        RECT 29.8 12 30.46 12.66 ;
      LAYER Metal4 ;
        RECT 29.8 12 30.46 12.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 270.44 12 271.1 12.66 ;
      LAYER Metal6 ;
        RECT 270.44 12 271.1 12.66 ;
      LAYER Metal3 ;
        RECT 270.44 12 271.1 12.66 ;
      LAYER Metal4 ;
        RECT 270.44 12 271.1 12.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 278.18 12 278.84 12.66 ;
      LAYER Metal6 ;
        RECT 278.18 12 278.84 12.66 ;
      LAYER Metal3 ;
        RECT 278.18 12 278.84 12.66 ;
      LAYER Metal4 ;
        RECT 278.18 12 278.84 12.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 291.72 12 292.38 12.66 ;
      LAYER Metal6 ;
        RECT 291.72 12 292.38 12.66 ;
      LAYER Metal3 ;
        RECT 291.72 12 292.38 12.66 ;
      LAYER Metal4 ;
        RECT 291.72 12 292.38 12.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 299.46 12 300.12 12.66 ;
      LAYER Metal6 ;
        RECT 299.46 12 300.12 12.66 ;
      LAYER Metal3 ;
        RECT 299.46 12 300.12 12.66 ;
      LAYER Metal4 ;
        RECT 299.46 12 300.12 12.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 313 12 313.66 12.66 ;
      LAYER Metal6 ;
        RECT 313 12 313.66 12.66 ;
      LAYER Metal3 ;
        RECT 313 12 313.66 12.66 ;
      LAYER Metal4 ;
        RECT 313 12 313.66 12.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 320.74 12 321.4 12.66 ;
      LAYER Metal6 ;
        RECT 320.74 12 321.4 12.66 ;
      LAYER Metal3 ;
        RECT 320.74 12 321.4 12.66 ;
      LAYER Metal4 ;
        RECT 320.74 12 321.4 12.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 334.28 12 334.94 12.66 ;
      LAYER Metal6 ;
        RECT 334.28 12 334.94 12.66 ;
      LAYER Metal3 ;
        RECT 334.28 12 334.94 12.66 ;
      LAYER Metal4 ;
        RECT 334.28 12 334.94 12.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 342.02 12 342.68 12.66 ;
      LAYER Metal6 ;
        RECT 342.02 12 342.68 12.66 ;
      LAYER Metal3 ;
        RECT 342.02 12 342.68 12.66 ;
      LAYER Metal4 ;
        RECT 342.02 12 342.68 12.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 355.56 12 356.22 12.66 ;
      LAYER Metal6 ;
        RECT 355.56 12 356.22 12.66 ;
      LAYER Metal3 ;
        RECT 355.56 12 356.22 12.66 ;
      LAYER Metal4 ;
        RECT 355.56 12 356.22 12.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 363.3 12 363.96 12.66 ;
      LAYER Metal6 ;
        RECT 363.3 12 363.96 12.66 ;
      LAYER Metal3 ;
        RECT 363.3 12 363.96 12.66 ;
      LAYER Metal4 ;
        RECT 363.3 12 363.96 12.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal6 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal3 ;
        RECT 43.34 12 44 12.66 ;
      LAYER Metal4 ;
        RECT 43.34 12 44 12.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 376.84 12 377.5 12.66 ;
      LAYER Metal6 ;
        RECT 376.84 12 377.5 12.66 ;
      LAYER Metal3 ;
        RECT 376.84 12 377.5 12.66 ;
      LAYER Metal4 ;
        RECT 376.84 12 377.5 12.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 384.58 12 385.24 12.66 ;
      LAYER Metal6 ;
        RECT 384.58 12 385.24 12.66 ;
      LAYER Metal3 ;
        RECT 384.58 12 385.24 12.66 ;
      LAYER Metal4 ;
        RECT 384.58 12 385.24 12.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal6 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal3 ;
        RECT 51.08 12 51.74 12.66 ;
      LAYER Metal4 ;
        RECT 51.08 12 51.74 12.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal6 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal3 ;
        RECT 64.62 12 65.28 12.66 ;
      LAYER Metal4 ;
        RECT 64.62 12 65.28 12.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal6 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal3 ;
        RECT 72.36 12 73.02 12.66 ;
      LAYER Metal4 ;
        RECT 72.36 12 73.02 12.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal6 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal3 ;
        RECT 85.9 12 86.56 12.66 ;
      LAYER Metal4 ;
        RECT 85.9 12 86.56 12.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal6 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal3 ;
        RECT 93.64 12 94.3 12.66 ;
      LAYER Metal4 ;
        RECT 93.64 12 94.3 12.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal6 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal3 ;
        RECT 107.18 12 107.84 12.66 ;
      LAYER Metal4 ;
        RECT 107.18 12 107.84 12.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal6 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal3 ;
        RECT 114.92 12 115.58 12.66 ;
      LAYER Metal4 ;
        RECT 114.92 12 115.58 12.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 212.68 12 213.34 12.66 ;
      LAYER Metal6 ;
        RECT 212.68 12 213.34 12.66 ;
      LAYER Metal3 ;
        RECT 212.68 12 213.34 12.66 ;
      LAYER Metal4 ;
        RECT 212.68 12 213.34 12.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal6 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal3 ;
        RECT 193.96 12 194.62 12.66 ;
      LAYER Metal4 ;
        RECT 193.96 12 194.62 12.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 140.035 423.015 145.035 ;
        RECT 0 0 423.015 5 ;
      LAYER Metal2 ;
        RECT 418.015 0 423.015 145.035 ;
        RECT 0 0 5 145.035 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 134.435 417.415 139.435 ;
        RECT 5.6 5.6 417.415 10.6 ;
      LAYER Metal2 ;
        RECT 412.415 5.6 417.415 139.435 ;
        RECT 5.6 5.6 10.6 139.435 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal2 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal3 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal4 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal5 ;
      RECT 12 12 411.02 132.965 ;
    LAYER Metal6 ;
      RECT 12 12 411.02 132.965 ;
  END
END MEM2_128X32

END LIBRARY
