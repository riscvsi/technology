VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;


MACRO MEM2_4096X32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM2_4096X32 0 0 ;
  SIZE 806.03 BY 947.445 ;
  SYMMETRY X Y R90 ;
  PIN A1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 287.155 13.46 287.815 ;
      LAYER Metal4 ;
        RECT 12.8 287.155 13.46 287.815 ;
      LAYER Metal5 ;
        RECT 12.8 287.155 13.46 287.815 ;
      LAYER Metal6 ;
        RECT 12.8 287.155 13.46 287.815 ;
    END
  END A1[0]
  PIN A1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 244.315 13.46 244.975 ;
      LAYER Metal4 ;
        RECT 12.8 244.315 13.46 244.975 ;
      LAYER Metal5 ;
        RECT 12.8 244.315 13.46 244.975 ;
      LAYER Metal6 ;
        RECT 12.8 244.315 13.46 244.975 ;
    END
  END A1[10]
  PIN A1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 241.215 13.46 241.875 ;
      LAYER Metal4 ;
        RECT 12.8 241.215 13.46 241.875 ;
      LAYER Metal5 ;
        RECT 12.8 241.215 13.46 241.875 ;
      LAYER Metal6 ;
        RECT 12.8 241.215 13.46 241.875 ;
    END
  END A1[11]
  PIN A1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 281.035 13.46 281.695 ;
      LAYER Metal4 ;
        RECT 12.8 281.035 13.46 281.695 ;
      LAYER Metal5 ;
        RECT 12.8 281.035 13.46 281.695 ;
      LAYER Metal6 ;
        RECT 12.8 281.035 13.46 281.695 ;
    END
  END A1[1]
  PIN A1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 277.935 13.46 278.595 ;
      LAYER Metal4 ;
        RECT 12.8 277.935 13.46 278.595 ;
      LAYER Metal5 ;
        RECT 12.8 277.935 13.46 278.595 ;
      LAYER Metal6 ;
        RECT 12.8 277.935 13.46 278.595 ;
    END
  END A1[2]
  PIN A1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 271.815 13.46 272.475 ;
      LAYER Metal4 ;
        RECT 12.8 271.815 13.46 272.475 ;
      LAYER Metal5 ;
        RECT 12.8 271.815 13.46 272.475 ;
      LAYER Metal6 ;
        RECT 12.8 271.815 13.46 272.475 ;
    END
  END A1[3]
  PIN A1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 268.795 13.46 269.455 ;
      LAYER Metal4 ;
        RECT 12.8 268.795 13.46 269.455 ;
      LAYER Metal5 ;
        RECT 12.8 268.795 13.46 269.455 ;
      LAYER Metal6 ;
        RECT 12.8 268.795 13.46 269.455 ;
    END
  END A1[4]
  PIN A1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 265.695 13.46 266.355 ;
      LAYER Metal4 ;
        RECT 12.8 265.695 13.46 266.355 ;
      LAYER Metal5 ;
        RECT 12.8 265.695 13.46 266.355 ;
      LAYER Metal6 ;
        RECT 12.8 265.695 13.46 266.355 ;
    END
  END A1[5]
  PIN A1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 259.575 13.46 260.235 ;
      LAYER Metal4 ;
        RECT 12.8 259.575 13.46 260.235 ;
      LAYER Metal5 ;
        RECT 12.8 259.575 13.46 260.235 ;
      LAYER Metal6 ;
        RECT 12.8 259.575 13.46 260.235 ;
    END
  END A1[6]
  PIN A1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 256.555 13.46 257.215 ;
      LAYER Metal4 ;
        RECT 12.8 256.555 13.46 257.215 ;
      LAYER Metal5 ;
        RECT 12.8 256.555 13.46 257.215 ;
      LAYER Metal6 ;
        RECT 12.8 256.555 13.46 257.215 ;
    END
  END A1[7]
  PIN A1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 253.455 13.46 254.115 ;
      LAYER Metal4 ;
        RECT 12.8 253.455 13.46 254.115 ;
      LAYER Metal5 ;
        RECT 12.8 253.455 13.46 254.115 ;
      LAYER Metal6 ;
        RECT 12.8 253.455 13.46 254.115 ;
    END
  END A1[8]
  PIN A1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 247.335 13.46 247.995 ;
      LAYER Metal4 ;
        RECT 12.8 247.335 13.46 247.995 ;
      LAYER Metal5 ;
        RECT 12.8 247.335 13.46 247.995 ;
      LAYER Metal6 ;
        RECT 12.8 247.335 13.46 247.995 ;
    END
  END A1[9]
  PIN A2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 111.515 13.46 112.175 ;
      LAYER Metal4 ;
        RECT 12.8 111.515 13.46 112.175 ;
      LAYER Metal5 ;
        RECT 12.8 111.515 13.46 112.175 ;
      LAYER Metal6 ;
        RECT 12.8 111.515 13.46 112.175 ;
    END
  END A2[0]
  PIN A2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 154.355 13.46 155.015 ;
      LAYER Metal4 ;
        RECT 12.8 154.355 13.46 155.015 ;
      LAYER Metal5 ;
        RECT 12.8 154.355 13.46 155.015 ;
      LAYER Metal6 ;
        RECT 12.8 154.355 13.46 155.015 ;
    END
  END A2[10]
  PIN A2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 157.455 13.46 158.115 ;
      LAYER Metal4 ;
        RECT 12.8 157.455 13.46 158.115 ;
      LAYER Metal5 ;
        RECT 12.8 157.455 13.46 158.115 ;
      LAYER Metal6 ;
        RECT 12.8 157.455 13.46 158.115 ;
    END
  END A2[11]
  PIN A2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 117.635 13.46 118.295 ;
      LAYER Metal4 ;
        RECT 12.8 117.635 13.46 118.295 ;
      LAYER Metal5 ;
        RECT 12.8 117.635 13.46 118.295 ;
      LAYER Metal6 ;
        RECT 12.8 117.635 13.46 118.295 ;
    END
  END A2[1]
  PIN A2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 120.735 13.46 121.395 ;
      LAYER Metal4 ;
        RECT 12.8 120.735 13.46 121.395 ;
      LAYER Metal5 ;
        RECT 12.8 120.735 13.46 121.395 ;
      LAYER Metal6 ;
        RECT 12.8 120.735 13.46 121.395 ;
    END
  END A2[2]
  PIN A2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 126.855 13.46 127.515 ;
      LAYER Metal4 ;
        RECT 12.8 126.855 13.46 127.515 ;
      LAYER Metal5 ;
        RECT 12.8 126.855 13.46 127.515 ;
      LAYER Metal6 ;
        RECT 12.8 126.855 13.46 127.515 ;
    END
  END A2[3]
  PIN A2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 129.875 13.46 130.535 ;
      LAYER Metal4 ;
        RECT 12.8 129.875 13.46 130.535 ;
      LAYER Metal5 ;
        RECT 12.8 129.875 13.46 130.535 ;
      LAYER Metal6 ;
        RECT 12.8 129.875 13.46 130.535 ;
    END
  END A2[4]
  PIN A2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 132.975 13.46 133.635 ;
      LAYER Metal4 ;
        RECT 12.8 132.975 13.46 133.635 ;
      LAYER Metal5 ;
        RECT 12.8 132.975 13.46 133.635 ;
      LAYER Metal6 ;
        RECT 12.8 132.975 13.46 133.635 ;
    END
  END A2[5]
  PIN A2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 139.095 13.46 139.755 ;
      LAYER Metal4 ;
        RECT 12.8 139.095 13.46 139.755 ;
      LAYER Metal5 ;
        RECT 12.8 139.095 13.46 139.755 ;
      LAYER Metal6 ;
        RECT 12.8 139.095 13.46 139.755 ;
    END
  END A2[6]
  PIN A2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 142.115 13.46 142.775 ;
      LAYER Metal4 ;
        RECT 12.8 142.115 13.46 142.775 ;
      LAYER Metal5 ;
        RECT 12.8 142.115 13.46 142.775 ;
      LAYER Metal6 ;
        RECT 12.8 142.115 13.46 142.775 ;
    END
  END A2[7]
  PIN A2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 145.215 13.46 145.875 ;
      LAYER Metal4 ;
        RECT 12.8 145.215 13.46 145.875 ;
      LAYER Metal5 ;
        RECT 12.8 145.215 13.46 145.875 ;
      LAYER Metal6 ;
        RECT 12.8 145.215 13.46 145.875 ;
    END
  END A2[8]
  PIN A2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 12.8 151.335 13.46 151.995 ;
      LAYER Metal4 ;
        RECT 12.8 151.335 13.46 151.995 ;
      LAYER Metal5 ;
        RECT 12.8 151.335 13.46 151.995 ;
      LAYER Metal6 ;
        RECT 12.8 151.335 13.46 151.995 ;
    END
  END A2[9]
  PIN CE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 395.57 13 396.23 13.66 ;
      LAYER Metal4 ;
        RECT 395.57 13 396.23 13.66 ;
      LAYER Metal5 ;
        RECT 395.57 13 396.23 13.66 ;
      LAYER Metal6 ;
        RECT 395.57 13 396.23 13.66 ;
    END
  END CE1
  PIN CE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 366.6 13 367.26 13.66 ;
      LAYER Metal4 ;
        RECT 366.6 13 367.26 13.66 ;
      LAYER Metal5 ;
        RECT 366.6 13 367.26 13.66 ;
      LAYER Metal6 ;
        RECT 366.6 13 367.26 13.66 ;
    END
  END CE2
  PIN CK1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 404.195 13 404.855 13.66 ;
      LAYER Metal4 ;
        RECT 404.195 13 404.855 13.66 ;
      LAYER Metal5 ;
        RECT 404.195 13 404.855 13.66 ;
      LAYER Metal6 ;
        RECT 404.195 13 404.855 13.66 ;
    END
  END CK1
  PIN CK2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 357.975 13 358.635 13.66 ;
      LAYER Metal4 ;
        RECT 357.975 13 358.635 13.66 ;
      LAYER Metal5 ;
        RECT 357.975 13 358.635 13.66 ;
      LAYER Metal6 ;
        RECT 357.975 13 358.635 13.66 ;
    END
  END CK2
  PIN D1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 21.91 13 22.57 13.66 ;
      LAYER Metal4 ;
        RECT 21.91 13 22.57 13.66 ;
      LAYER Metal5 ;
        RECT 21.91 13 22.57 13.66 ;
      LAYER Metal6 ;
        RECT 21.91 13 22.57 13.66 ;
    END
  END D1[0]
  PIN D1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 234.71 13 235.37 13.66 ;
      LAYER Metal4 ;
        RECT 234.71 13 235.37 13.66 ;
      LAYER Metal5 ;
        RECT 234.71 13 235.37 13.66 ;
      LAYER Metal6 ;
        RECT 234.71 13 235.37 13.66 ;
    END
  END D1[10]
  PIN D1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 264.03 13 264.69 13.66 ;
      LAYER Metal4 ;
        RECT 264.03 13 264.69 13.66 ;
      LAYER Metal5 ;
        RECT 264.03 13 264.69 13.66 ;
      LAYER Metal6 ;
        RECT 264.03 13 264.69 13.66 ;
    END
  END D1[11]
  PIN D1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 277.27 13 277.93 13.66 ;
      LAYER Metal4 ;
        RECT 277.27 13 277.93 13.66 ;
      LAYER Metal5 ;
        RECT 277.27 13 277.93 13.66 ;
      LAYER Metal6 ;
        RECT 277.27 13 277.93 13.66 ;
    END
  END D1[12]
  PIN D1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 306.59 13 307.25 13.66 ;
      LAYER Metal4 ;
        RECT 306.59 13 307.25 13.66 ;
      LAYER Metal5 ;
        RECT 306.59 13 307.25 13.66 ;
      LAYER Metal6 ;
        RECT 306.59 13 307.25 13.66 ;
    END
  END D1[13]
  PIN D1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 319.83 13 320.49 13.66 ;
      LAYER Metal4 ;
        RECT 319.83 13 320.49 13.66 ;
      LAYER Metal5 ;
        RECT 319.83 13 320.49 13.66 ;
      LAYER Metal6 ;
        RECT 319.83 13 320.49 13.66 ;
    END
  END D1[14]
  PIN D1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 349.15 13 349.81 13.66 ;
      LAYER Metal4 ;
        RECT 349.15 13 349.81 13.66 ;
      LAYER Metal5 ;
        RECT 349.15 13 349.81 13.66 ;
      LAYER Metal6 ;
        RECT 349.15 13 349.81 13.66 ;
    END
  END D1[15]
  PIN D1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 413.02 13 413.68 13.66 ;
      LAYER Metal4 ;
        RECT 413.02 13 413.68 13.66 ;
      LAYER Metal5 ;
        RECT 413.02 13 413.68 13.66 ;
      LAYER Metal6 ;
        RECT 413.02 13 413.68 13.66 ;
    END
  END D1[16]
  PIN D1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 442.34 13 443 13.66 ;
      LAYER Metal4 ;
        RECT 442.34 13 443 13.66 ;
      LAYER Metal5 ;
        RECT 442.34 13 443 13.66 ;
      LAYER Metal6 ;
        RECT 442.34 13 443 13.66 ;
    END
  END D1[17]
  PIN D1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 455.58 13 456.24 13.66 ;
      LAYER Metal4 ;
        RECT 455.58 13 456.24 13.66 ;
      LAYER Metal5 ;
        RECT 455.58 13 456.24 13.66 ;
      LAYER Metal6 ;
        RECT 455.58 13 456.24 13.66 ;
    END
  END D1[18]
  PIN D1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 484.9 13 485.56 13.66 ;
      LAYER Metal4 ;
        RECT 484.9 13 485.56 13.66 ;
      LAYER Metal5 ;
        RECT 484.9 13 485.56 13.66 ;
      LAYER Metal6 ;
        RECT 484.9 13 485.56 13.66 ;
    END
  END D1[19]
  PIN D1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 51.23 13 51.89 13.66 ;
      LAYER Metal4 ;
        RECT 51.23 13 51.89 13.66 ;
      LAYER Metal5 ;
        RECT 51.23 13 51.89 13.66 ;
      LAYER Metal6 ;
        RECT 51.23 13 51.89 13.66 ;
    END
  END D1[1]
  PIN D1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 498.14 13 498.8 13.66 ;
      LAYER Metal4 ;
        RECT 498.14 13 498.8 13.66 ;
      LAYER Metal5 ;
        RECT 498.14 13 498.8 13.66 ;
      LAYER Metal6 ;
        RECT 498.14 13 498.8 13.66 ;
    END
  END D1[20]
  PIN D1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 527.46 13 528.12 13.66 ;
      LAYER Metal4 ;
        RECT 527.46 13 528.12 13.66 ;
      LAYER Metal5 ;
        RECT 527.46 13 528.12 13.66 ;
      LAYER Metal6 ;
        RECT 527.46 13 528.12 13.66 ;
    END
  END D1[21]
  PIN D1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 540.7 13 541.36 13.66 ;
      LAYER Metal4 ;
        RECT 540.7 13 541.36 13.66 ;
      LAYER Metal5 ;
        RECT 540.7 13 541.36 13.66 ;
      LAYER Metal6 ;
        RECT 540.7 13 541.36 13.66 ;
    END
  END D1[22]
  PIN D1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 570.02 13 570.68 13.66 ;
      LAYER Metal4 ;
        RECT 570.02 13 570.68 13.66 ;
      LAYER Metal5 ;
        RECT 570.02 13 570.68 13.66 ;
      LAYER Metal6 ;
        RECT 570.02 13 570.68 13.66 ;
    END
  END D1[23]
  PIN D1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 583.26 13 583.92 13.66 ;
      LAYER Metal4 ;
        RECT 583.26 13 583.92 13.66 ;
      LAYER Metal5 ;
        RECT 583.26 13 583.92 13.66 ;
      LAYER Metal6 ;
        RECT 583.26 13 583.92 13.66 ;
    END
  END D1[24]
  PIN D1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 612.58 13 613.24 13.66 ;
      LAYER Metal4 ;
        RECT 612.58 13 613.24 13.66 ;
      LAYER Metal5 ;
        RECT 612.58 13 613.24 13.66 ;
      LAYER Metal6 ;
        RECT 612.58 13 613.24 13.66 ;
    END
  END D1[25]
  PIN D1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 625.82 13 626.48 13.66 ;
      LAYER Metal4 ;
        RECT 625.82 13 626.48 13.66 ;
      LAYER Metal5 ;
        RECT 625.82 13 626.48 13.66 ;
      LAYER Metal6 ;
        RECT 625.82 13 626.48 13.66 ;
    END
  END D1[26]
  PIN D1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 655.14 13 655.8 13.66 ;
      LAYER Metal4 ;
        RECT 655.14 13 655.8 13.66 ;
      LAYER Metal5 ;
        RECT 655.14 13 655.8 13.66 ;
      LAYER Metal6 ;
        RECT 655.14 13 655.8 13.66 ;
    END
  END D1[27]
  PIN D1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 668.38 13 669.04 13.66 ;
      LAYER Metal4 ;
        RECT 668.38 13 669.04 13.66 ;
      LAYER Metal5 ;
        RECT 668.38 13 669.04 13.66 ;
      LAYER Metal6 ;
        RECT 668.38 13 669.04 13.66 ;
    END
  END D1[28]
  PIN D1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 697.7 13 698.36 13.66 ;
      LAYER Metal4 ;
        RECT 697.7 13 698.36 13.66 ;
      LAYER Metal5 ;
        RECT 697.7 13 698.36 13.66 ;
      LAYER Metal6 ;
        RECT 697.7 13 698.36 13.66 ;
    END
  END D1[29]
  PIN D1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 64.47 13 65.13 13.66 ;
      LAYER Metal4 ;
        RECT 64.47 13 65.13 13.66 ;
      LAYER Metal5 ;
        RECT 64.47 13 65.13 13.66 ;
      LAYER Metal6 ;
        RECT 64.47 13 65.13 13.66 ;
    END
  END D1[2]
  PIN D1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 710.94 13 711.6 13.66 ;
      LAYER Metal4 ;
        RECT 710.94 13 711.6 13.66 ;
      LAYER Metal5 ;
        RECT 710.94 13 711.6 13.66 ;
      LAYER Metal6 ;
        RECT 710.94 13 711.6 13.66 ;
    END
  END D1[30]
  PIN D1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 740.26 13 740.92 13.66 ;
      LAYER Metal4 ;
        RECT 740.26 13 740.92 13.66 ;
      LAYER Metal5 ;
        RECT 740.26 13 740.92 13.66 ;
      LAYER Metal6 ;
        RECT 740.26 13 740.92 13.66 ;
    END
  END D1[31]
  PIN D1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 93.79 13 94.45 13.66 ;
      LAYER Metal4 ;
        RECT 93.79 13 94.45 13.66 ;
      LAYER Metal5 ;
        RECT 93.79 13 94.45 13.66 ;
      LAYER Metal6 ;
        RECT 93.79 13 94.45 13.66 ;
    END
  END D1[3]
  PIN D1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 107.03 13 107.69 13.66 ;
      LAYER Metal4 ;
        RECT 107.03 13 107.69 13.66 ;
      LAYER Metal5 ;
        RECT 107.03 13 107.69 13.66 ;
      LAYER Metal6 ;
        RECT 107.03 13 107.69 13.66 ;
    END
  END D1[4]
  PIN D1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 136.35 13 137.01 13.66 ;
      LAYER Metal4 ;
        RECT 136.35 13 137.01 13.66 ;
      LAYER Metal5 ;
        RECT 136.35 13 137.01 13.66 ;
      LAYER Metal6 ;
        RECT 136.35 13 137.01 13.66 ;
    END
  END D1[5]
  PIN D1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 149.59 13 150.25 13.66 ;
      LAYER Metal4 ;
        RECT 149.59 13 150.25 13.66 ;
      LAYER Metal5 ;
        RECT 149.59 13 150.25 13.66 ;
      LAYER Metal6 ;
        RECT 149.59 13 150.25 13.66 ;
    END
  END D1[6]
  PIN D1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 178.91 13 179.57 13.66 ;
      LAYER Metal4 ;
        RECT 178.91 13 179.57 13.66 ;
      LAYER Metal5 ;
        RECT 178.91 13 179.57 13.66 ;
      LAYER Metal6 ;
        RECT 178.91 13 179.57 13.66 ;
    END
  END D1[7]
  PIN D1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 192.15 13 192.81 13.66 ;
      LAYER Metal4 ;
        RECT 192.15 13 192.81 13.66 ;
      LAYER Metal5 ;
        RECT 192.15 13 192.81 13.66 ;
      LAYER Metal6 ;
        RECT 192.15 13 192.81 13.66 ;
    END
  END D1[8]
  PIN D1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 221.47 13 222.13 13.66 ;
      LAYER Metal4 ;
        RECT 221.47 13 222.13 13.66 ;
      LAYER Metal5 ;
        RECT 221.47 13 222.13 13.66 ;
      LAYER Metal6 ;
        RECT 221.47 13 222.13 13.66 ;
    END
  END D1[9]
  PIN D2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 29.95 13 30.61 13.66 ;
      LAYER Metal4 ;
        RECT 29.95 13 30.61 13.66 ;
      LAYER Metal5 ;
        RECT 29.95 13 30.61 13.66 ;
      LAYER Metal6 ;
        RECT 29.95 13 30.61 13.66 ;
    END
  END D2[0]
  PIN D2[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 242.75 13 243.41 13.66 ;
      LAYER Metal4 ;
        RECT 242.75 13 243.41 13.66 ;
      LAYER Metal5 ;
        RECT 242.75 13 243.41 13.66 ;
      LAYER Metal6 ;
        RECT 242.75 13 243.41 13.66 ;
    END
  END D2[10]
  PIN D2[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 255.99 13 256.65 13.66 ;
      LAYER Metal4 ;
        RECT 255.99 13 256.65 13.66 ;
      LAYER Metal5 ;
        RECT 255.99 13 256.65 13.66 ;
      LAYER Metal6 ;
        RECT 255.99 13 256.65 13.66 ;
    END
  END D2[11]
  PIN D2[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 285.31 13 285.97 13.66 ;
      LAYER Metal4 ;
        RECT 285.31 13 285.97 13.66 ;
      LAYER Metal5 ;
        RECT 285.31 13 285.97 13.66 ;
      LAYER Metal6 ;
        RECT 285.31 13 285.97 13.66 ;
    END
  END D2[12]
  PIN D2[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 298.55 13 299.21 13.66 ;
      LAYER Metal4 ;
        RECT 298.55 13 299.21 13.66 ;
      LAYER Metal5 ;
        RECT 298.55 13 299.21 13.66 ;
      LAYER Metal6 ;
        RECT 298.55 13 299.21 13.66 ;
    END
  END D2[13]
  PIN D2[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 327.87 13 328.53 13.66 ;
      LAYER Metal4 ;
        RECT 327.87 13 328.53 13.66 ;
      LAYER Metal5 ;
        RECT 327.87 13 328.53 13.66 ;
      LAYER Metal6 ;
        RECT 327.87 13 328.53 13.66 ;
    END
  END D2[14]
  PIN D2[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 341.11 13 341.77 13.66 ;
      LAYER Metal4 ;
        RECT 341.11 13 341.77 13.66 ;
      LAYER Metal5 ;
        RECT 341.11 13 341.77 13.66 ;
      LAYER Metal6 ;
        RECT 341.11 13 341.77 13.66 ;
    END
  END D2[15]
  PIN D2[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 421.06 13 421.72 13.66 ;
      LAYER Metal4 ;
        RECT 421.06 13 421.72 13.66 ;
      LAYER Metal5 ;
        RECT 421.06 13 421.72 13.66 ;
      LAYER Metal6 ;
        RECT 421.06 13 421.72 13.66 ;
    END
  END D2[16]
  PIN D2[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 434.3 13 434.96 13.66 ;
      LAYER Metal4 ;
        RECT 434.3 13 434.96 13.66 ;
      LAYER Metal5 ;
        RECT 434.3 13 434.96 13.66 ;
      LAYER Metal6 ;
        RECT 434.3 13 434.96 13.66 ;
    END
  END D2[17]
  PIN D2[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 463.62 13 464.28 13.66 ;
      LAYER Metal4 ;
        RECT 463.62 13 464.28 13.66 ;
      LAYER Metal5 ;
        RECT 463.62 13 464.28 13.66 ;
      LAYER Metal6 ;
        RECT 463.62 13 464.28 13.66 ;
    END
  END D2[18]
  PIN D2[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 476.86 13 477.52 13.66 ;
      LAYER Metal4 ;
        RECT 476.86 13 477.52 13.66 ;
      LAYER Metal5 ;
        RECT 476.86 13 477.52 13.66 ;
      LAYER Metal6 ;
        RECT 476.86 13 477.52 13.66 ;
    END
  END D2[19]
  PIN D2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 43.19 13 43.85 13.66 ;
      LAYER Metal4 ;
        RECT 43.19 13 43.85 13.66 ;
      LAYER Metal5 ;
        RECT 43.19 13 43.85 13.66 ;
      LAYER Metal6 ;
        RECT 43.19 13 43.85 13.66 ;
    END
  END D2[1]
  PIN D2[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 506.18 13 506.84 13.66 ;
      LAYER Metal4 ;
        RECT 506.18 13 506.84 13.66 ;
      LAYER Metal5 ;
        RECT 506.18 13 506.84 13.66 ;
      LAYER Metal6 ;
        RECT 506.18 13 506.84 13.66 ;
    END
  END D2[20]
  PIN D2[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 519.42 13 520.08 13.66 ;
      LAYER Metal4 ;
        RECT 519.42 13 520.08 13.66 ;
      LAYER Metal5 ;
        RECT 519.42 13 520.08 13.66 ;
      LAYER Metal6 ;
        RECT 519.42 13 520.08 13.66 ;
    END
  END D2[21]
  PIN D2[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 548.74 13 549.4 13.66 ;
      LAYER Metal4 ;
        RECT 548.74 13 549.4 13.66 ;
      LAYER Metal5 ;
        RECT 548.74 13 549.4 13.66 ;
      LAYER Metal6 ;
        RECT 548.74 13 549.4 13.66 ;
    END
  END D2[22]
  PIN D2[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 561.98 13 562.64 13.66 ;
      LAYER Metal4 ;
        RECT 561.98 13 562.64 13.66 ;
      LAYER Metal5 ;
        RECT 561.98 13 562.64 13.66 ;
      LAYER Metal6 ;
        RECT 561.98 13 562.64 13.66 ;
    END
  END D2[23]
  PIN D2[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 591.3 13 591.96 13.66 ;
      LAYER Metal4 ;
        RECT 591.3 13 591.96 13.66 ;
      LAYER Metal5 ;
        RECT 591.3 13 591.96 13.66 ;
      LAYER Metal6 ;
        RECT 591.3 13 591.96 13.66 ;
    END
  END D2[24]
  PIN D2[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 604.54 13 605.2 13.66 ;
      LAYER Metal4 ;
        RECT 604.54 13 605.2 13.66 ;
      LAYER Metal5 ;
        RECT 604.54 13 605.2 13.66 ;
      LAYER Metal6 ;
        RECT 604.54 13 605.2 13.66 ;
    END
  END D2[25]
  PIN D2[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 633.86 13 634.52 13.66 ;
      LAYER Metal4 ;
        RECT 633.86 13 634.52 13.66 ;
      LAYER Metal5 ;
        RECT 633.86 13 634.52 13.66 ;
      LAYER Metal6 ;
        RECT 633.86 13 634.52 13.66 ;
    END
  END D2[26]
  PIN D2[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 647.1 13 647.76 13.66 ;
      LAYER Metal4 ;
        RECT 647.1 13 647.76 13.66 ;
      LAYER Metal5 ;
        RECT 647.1 13 647.76 13.66 ;
      LAYER Metal6 ;
        RECT 647.1 13 647.76 13.66 ;
    END
  END D2[27]
  PIN D2[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 676.42 13 677.08 13.66 ;
      LAYER Metal4 ;
        RECT 676.42 13 677.08 13.66 ;
      LAYER Metal5 ;
        RECT 676.42 13 677.08 13.66 ;
      LAYER Metal6 ;
        RECT 676.42 13 677.08 13.66 ;
    END
  END D2[28]
  PIN D2[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 689.66 13 690.32 13.66 ;
      LAYER Metal4 ;
        RECT 689.66 13 690.32 13.66 ;
      LAYER Metal5 ;
        RECT 689.66 13 690.32 13.66 ;
      LAYER Metal6 ;
        RECT 689.66 13 690.32 13.66 ;
    END
  END D2[29]
  PIN D2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 72.51 13 73.17 13.66 ;
      LAYER Metal4 ;
        RECT 72.51 13 73.17 13.66 ;
      LAYER Metal5 ;
        RECT 72.51 13 73.17 13.66 ;
      LAYER Metal6 ;
        RECT 72.51 13 73.17 13.66 ;
    END
  END D2[2]
  PIN D2[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 718.98 13 719.64 13.66 ;
      LAYER Metal4 ;
        RECT 718.98 13 719.64 13.66 ;
      LAYER Metal5 ;
        RECT 718.98 13 719.64 13.66 ;
      LAYER Metal6 ;
        RECT 718.98 13 719.64 13.66 ;
    END
  END D2[30]
  PIN D2[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 732.22 13 732.88 13.66 ;
      LAYER Metal4 ;
        RECT 732.22 13 732.88 13.66 ;
      LAYER Metal5 ;
        RECT 732.22 13 732.88 13.66 ;
      LAYER Metal6 ;
        RECT 732.22 13 732.88 13.66 ;
    END
  END D2[31]
  PIN D2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 85.75 13 86.41 13.66 ;
      LAYER Metal4 ;
        RECT 85.75 13 86.41 13.66 ;
      LAYER Metal5 ;
        RECT 85.75 13 86.41 13.66 ;
      LAYER Metal6 ;
        RECT 85.75 13 86.41 13.66 ;
    END
  END D2[3]
  PIN D2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 115.07 13 115.73 13.66 ;
      LAYER Metal4 ;
        RECT 115.07 13 115.73 13.66 ;
      LAYER Metal5 ;
        RECT 115.07 13 115.73 13.66 ;
      LAYER Metal6 ;
        RECT 115.07 13 115.73 13.66 ;
    END
  END D2[4]
  PIN D2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 128.31 13 128.97 13.66 ;
      LAYER Metal4 ;
        RECT 128.31 13 128.97 13.66 ;
      LAYER Metal5 ;
        RECT 128.31 13 128.97 13.66 ;
      LAYER Metal6 ;
        RECT 128.31 13 128.97 13.66 ;
    END
  END D2[5]
  PIN D2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 157.63 13 158.29 13.66 ;
      LAYER Metal4 ;
        RECT 157.63 13 158.29 13.66 ;
      LAYER Metal5 ;
        RECT 157.63 13 158.29 13.66 ;
      LAYER Metal6 ;
        RECT 157.63 13 158.29 13.66 ;
    END
  END D2[6]
  PIN D2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 170.87 13 171.53 13.66 ;
      LAYER Metal4 ;
        RECT 170.87 13 171.53 13.66 ;
      LAYER Metal5 ;
        RECT 170.87 13 171.53 13.66 ;
      LAYER Metal6 ;
        RECT 170.87 13 171.53 13.66 ;
    END
  END D2[7]
  PIN D2[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 200.19 13 200.85 13.66 ;
      LAYER Metal4 ;
        RECT 200.19 13 200.85 13.66 ;
      LAYER Metal5 ;
        RECT 200.19 13 200.85 13.66 ;
      LAYER Metal6 ;
        RECT 200.19 13 200.85 13.66 ;
    END
  END D2[8]
  PIN D2[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 213.43 13 214.09 13.66 ;
      LAYER Metal4 ;
        RECT 213.43 13 214.09 13.66 ;
      LAYER Metal5 ;
        RECT 213.43 13 214.09 13.66 ;
      LAYER Metal6 ;
        RECT 213.43 13 214.09 13.66 ;
    END
  END D2[9]
  PIN Q1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 24.49 13 25.15 13.66 ;
      LAYER Metal4 ;
        RECT 24.49 13 25.15 13.66 ;
      LAYER Metal5 ;
        RECT 24.49 13 25.15 13.66 ;
      LAYER Metal6 ;
        RECT 24.49 13 25.15 13.66 ;
    END
  END Q1[0]
  PIN Q1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 237.29 13 237.95 13.66 ;
      LAYER Metal4 ;
        RECT 237.29 13 237.95 13.66 ;
      LAYER Metal5 ;
        RECT 237.29 13 237.95 13.66 ;
      LAYER Metal6 ;
        RECT 237.29 13 237.95 13.66 ;
    END
  END Q1[10]
  PIN Q1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 261.45 13 262.11 13.66 ;
      LAYER Metal4 ;
        RECT 261.45 13 262.11 13.66 ;
      LAYER Metal5 ;
        RECT 261.45 13 262.11 13.66 ;
      LAYER Metal6 ;
        RECT 261.45 13 262.11 13.66 ;
    END
  END Q1[11]
  PIN Q1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 279.85 13 280.51 13.66 ;
      LAYER Metal4 ;
        RECT 279.85 13 280.51 13.66 ;
      LAYER Metal5 ;
        RECT 279.85 13 280.51 13.66 ;
      LAYER Metal6 ;
        RECT 279.85 13 280.51 13.66 ;
    END
  END Q1[12]
  PIN Q1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 304.01 13 304.67 13.66 ;
      LAYER Metal4 ;
        RECT 304.01 13 304.67 13.66 ;
      LAYER Metal5 ;
        RECT 304.01 13 304.67 13.66 ;
      LAYER Metal6 ;
        RECT 304.01 13 304.67 13.66 ;
    END
  END Q1[13]
  PIN Q1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 322.41 13 323.07 13.66 ;
      LAYER Metal4 ;
        RECT 322.41 13 323.07 13.66 ;
      LAYER Metal5 ;
        RECT 322.41 13 323.07 13.66 ;
      LAYER Metal6 ;
        RECT 322.41 13 323.07 13.66 ;
    END
  END Q1[14]
  PIN Q1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 346.57 13 347.23 13.66 ;
      LAYER Metal4 ;
        RECT 346.57 13 347.23 13.66 ;
      LAYER Metal5 ;
        RECT 346.57 13 347.23 13.66 ;
      LAYER Metal6 ;
        RECT 346.57 13 347.23 13.66 ;
    END
  END Q1[15]
  PIN Q1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 415.6 13 416.26 13.66 ;
      LAYER Metal4 ;
        RECT 415.6 13 416.26 13.66 ;
      LAYER Metal5 ;
        RECT 415.6 13 416.26 13.66 ;
      LAYER Metal6 ;
        RECT 415.6 13 416.26 13.66 ;
    END
  END Q1[16]
  PIN Q1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 439.76 13 440.42 13.66 ;
      LAYER Metal4 ;
        RECT 439.76 13 440.42 13.66 ;
      LAYER Metal5 ;
        RECT 439.76 13 440.42 13.66 ;
      LAYER Metal6 ;
        RECT 439.76 13 440.42 13.66 ;
    END
  END Q1[17]
  PIN Q1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 458.16 13 458.82 13.66 ;
      LAYER Metal4 ;
        RECT 458.16 13 458.82 13.66 ;
      LAYER Metal5 ;
        RECT 458.16 13 458.82 13.66 ;
      LAYER Metal6 ;
        RECT 458.16 13 458.82 13.66 ;
    END
  END Q1[18]
  PIN Q1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 482.32 13 482.98 13.66 ;
      LAYER Metal4 ;
        RECT 482.32 13 482.98 13.66 ;
      LAYER Metal5 ;
        RECT 482.32 13 482.98 13.66 ;
      LAYER Metal6 ;
        RECT 482.32 13 482.98 13.66 ;
    END
  END Q1[19]
  PIN Q1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 48.65 13 49.31 13.66 ;
      LAYER Metal4 ;
        RECT 48.65 13 49.31 13.66 ;
      LAYER Metal5 ;
        RECT 48.65 13 49.31 13.66 ;
      LAYER Metal6 ;
        RECT 48.65 13 49.31 13.66 ;
    END
  END Q1[1]
  PIN Q1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 500.72 13 501.38 13.66 ;
      LAYER Metal4 ;
        RECT 500.72 13 501.38 13.66 ;
      LAYER Metal5 ;
        RECT 500.72 13 501.38 13.66 ;
      LAYER Metal6 ;
        RECT 500.72 13 501.38 13.66 ;
    END
  END Q1[20]
  PIN Q1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 524.88 13 525.54 13.66 ;
      LAYER Metal4 ;
        RECT 524.88 13 525.54 13.66 ;
      LAYER Metal5 ;
        RECT 524.88 13 525.54 13.66 ;
      LAYER Metal6 ;
        RECT 524.88 13 525.54 13.66 ;
    END
  END Q1[21]
  PIN Q1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 543.28 13 543.94 13.66 ;
      LAYER Metal4 ;
        RECT 543.28 13 543.94 13.66 ;
      LAYER Metal5 ;
        RECT 543.28 13 543.94 13.66 ;
      LAYER Metal6 ;
        RECT 543.28 13 543.94 13.66 ;
    END
  END Q1[22]
  PIN Q1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 567.44 13 568.1 13.66 ;
      LAYER Metal4 ;
        RECT 567.44 13 568.1 13.66 ;
      LAYER Metal5 ;
        RECT 567.44 13 568.1 13.66 ;
      LAYER Metal6 ;
        RECT 567.44 13 568.1 13.66 ;
    END
  END Q1[23]
  PIN Q1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 585.84 13 586.5 13.66 ;
      LAYER Metal4 ;
        RECT 585.84 13 586.5 13.66 ;
      LAYER Metal5 ;
        RECT 585.84 13 586.5 13.66 ;
      LAYER Metal6 ;
        RECT 585.84 13 586.5 13.66 ;
    END
  END Q1[24]
  PIN Q1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 610 13 610.66 13.66 ;
      LAYER Metal4 ;
        RECT 610 13 610.66 13.66 ;
      LAYER Metal5 ;
        RECT 610 13 610.66 13.66 ;
      LAYER Metal6 ;
        RECT 610 13 610.66 13.66 ;
    END
  END Q1[25]
  PIN Q1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 628.4 13 629.06 13.66 ;
      LAYER Metal4 ;
        RECT 628.4 13 629.06 13.66 ;
      LAYER Metal5 ;
        RECT 628.4 13 629.06 13.66 ;
      LAYER Metal6 ;
        RECT 628.4 13 629.06 13.66 ;
    END
  END Q1[26]
  PIN Q1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 652.56 13 653.22 13.66 ;
      LAYER Metal4 ;
        RECT 652.56 13 653.22 13.66 ;
      LAYER Metal5 ;
        RECT 652.56 13 653.22 13.66 ;
      LAYER Metal6 ;
        RECT 652.56 13 653.22 13.66 ;
    END
  END Q1[27]
  PIN Q1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 670.96 13 671.62 13.66 ;
      LAYER Metal4 ;
        RECT 670.96 13 671.62 13.66 ;
      LAYER Metal5 ;
        RECT 670.96 13 671.62 13.66 ;
      LAYER Metal6 ;
        RECT 670.96 13 671.62 13.66 ;
    END
  END Q1[28]
  PIN Q1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 695.12 13 695.78 13.66 ;
      LAYER Metal4 ;
        RECT 695.12 13 695.78 13.66 ;
      LAYER Metal5 ;
        RECT 695.12 13 695.78 13.66 ;
      LAYER Metal6 ;
        RECT 695.12 13 695.78 13.66 ;
    END
  END Q1[29]
  PIN Q1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 67.05 13 67.71 13.66 ;
      LAYER Metal4 ;
        RECT 67.05 13 67.71 13.66 ;
      LAYER Metal5 ;
        RECT 67.05 13 67.71 13.66 ;
      LAYER Metal6 ;
        RECT 67.05 13 67.71 13.66 ;
    END
  END Q1[2]
  PIN Q1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 713.52 13 714.18 13.66 ;
      LAYER Metal4 ;
        RECT 713.52 13 714.18 13.66 ;
      LAYER Metal5 ;
        RECT 713.52 13 714.18 13.66 ;
      LAYER Metal6 ;
        RECT 713.52 13 714.18 13.66 ;
    END
  END Q1[30]
  PIN Q1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 737.68 13 738.34 13.66 ;
      LAYER Metal4 ;
        RECT 737.68 13 738.34 13.66 ;
      LAYER Metal5 ;
        RECT 737.68 13 738.34 13.66 ;
      LAYER Metal6 ;
        RECT 737.68 13 738.34 13.66 ;
    END
  END Q1[31]
  PIN Q1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 91.21 13 91.87 13.66 ;
      LAYER Metal4 ;
        RECT 91.21 13 91.87 13.66 ;
      LAYER Metal5 ;
        RECT 91.21 13 91.87 13.66 ;
      LAYER Metal6 ;
        RECT 91.21 13 91.87 13.66 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 109.61 13 110.27 13.66 ;
      LAYER Metal4 ;
        RECT 109.61 13 110.27 13.66 ;
      LAYER Metal5 ;
        RECT 109.61 13 110.27 13.66 ;
      LAYER Metal6 ;
        RECT 109.61 13 110.27 13.66 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 133.77 13 134.43 13.66 ;
      LAYER Metal4 ;
        RECT 133.77 13 134.43 13.66 ;
      LAYER Metal5 ;
        RECT 133.77 13 134.43 13.66 ;
      LAYER Metal6 ;
        RECT 133.77 13 134.43 13.66 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 152.17 13 152.83 13.66 ;
      LAYER Metal4 ;
        RECT 152.17 13 152.83 13.66 ;
      LAYER Metal5 ;
        RECT 152.17 13 152.83 13.66 ;
      LAYER Metal6 ;
        RECT 152.17 13 152.83 13.66 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 176.33 13 176.99 13.66 ;
      LAYER Metal4 ;
        RECT 176.33 13 176.99 13.66 ;
      LAYER Metal5 ;
        RECT 176.33 13 176.99 13.66 ;
      LAYER Metal6 ;
        RECT 176.33 13 176.99 13.66 ;
    END
  END Q1[7]
  PIN Q1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 194.73 13 195.39 13.66 ;
      LAYER Metal4 ;
        RECT 194.73 13 195.39 13.66 ;
      LAYER Metal5 ;
        RECT 194.73 13 195.39 13.66 ;
      LAYER Metal6 ;
        RECT 194.73 13 195.39 13.66 ;
    END
  END Q1[8]
  PIN Q1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 218.89 13 219.55 13.66 ;
      LAYER Metal4 ;
        RECT 218.89 13 219.55 13.66 ;
      LAYER Metal5 ;
        RECT 218.89 13 219.55 13.66 ;
      LAYER Metal6 ;
        RECT 218.89 13 219.55 13.66 ;
    END
  END Q1[9]
  PIN Q2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 27.37 13 28.03 13.66 ;
      LAYER Metal4 ;
        RECT 27.37 13 28.03 13.66 ;
      LAYER Metal5 ;
        RECT 27.37 13 28.03 13.66 ;
      LAYER Metal6 ;
        RECT 27.37 13 28.03 13.66 ;
    END
  END Q2[0]
  PIN Q2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 240.17 13 240.83 13.66 ;
      LAYER Metal4 ;
        RECT 240.17 13 240.83 13.66 ;
      LAYER Metal5 ;
        RECT 240.17 13 240.83 13.66 ;
      LAYER Metal6 ;
        RECT 240.17 13 240.83 13.66 ;
    END
  END Q2[10]
  PIN Q2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 258.57 13 259.23 13.66 ;
      LAYER Metal4 ;
        RECT 258.57 13 259.23 13.66 ;
      LAYER Metal5 ;
        RECT 258.57 13 259.23 13.66 ;
      LAYER Metal6 ;
        RECT 258.57 13 259.23 13.66 ;
    END
  END Q2[11]
  PIN Q2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 282.73 13 283.39 13.66 ;
      LAYER Metal4 ;
        RECT 282.73 13 283.39 13.66 ;
      LAYER Metal5 ;
        RECT 282.73 13 283.39 13.66 ;
      LAYER Metal6 ;
        RECT 282.73 13 283.39 13.66 ;
    END
  END Q2[12]
  PIN Q2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 301.13 13 301.79 13.66 ;
      LAYER Metal4 ;
        RECT 301.13 13 301.79 13.66 ;
      LAYER Metal5 ;
        RECT 301.13 13 301.79 13.66 ;
      LAYER Metal6 ;
        RECT 301.13 13 301.79 13.66 ;
    END
  END Q2[13]
  PIN Q2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 325.29 13 325.95 13.66 ;
      LAYER Metal4 ;
        RECT 325.29 13 325.95 13.66 ;
      LAYER Metal5 ;
        RECT 325.29 13 325.95 13.66 ;
      LAYER Metal6 ;
        RECT 325.29 13 325.95 13.66 ;
    END
  END Q2[14]
  PIN Q2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 343.69 13 344.35 13.66 ;
      LAYER Metal4 ;
        RECT 343.69 13 344.35 13.66 ;
      LAYER Metal5 ;
        RECT 343.69 13 344.35 13.66 ;
      LAYER Metal6 ;
        RECT 343.69 13 344.35 13.66 ;
    END
  END Q2[15]
  PIN Q2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 418.48 13 419.14 13.66 ;
      LAYER Metal4 ;
        RECT 418.48 13 419.14 13.66 ;
      LAYER Metal5 ;
        RECT 418.48 13 419.14 13.66 ;
      LAYER Metal6 ;
        RECT 418.48 13 419.14 13.66 ;
    END
  END Q2[16]
  PIN Q2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 436.88 13 437.54 13.66 ;
      LAYER Metal4 ;
        RECT 436.88 13 437.54 13.66 ;
      LAYER Metal5 ;
        RECT 436.88 13 437.54 13.66 ;
      LAYER Metal6 ;
        RECT 436.88 13 437.54 13.66 ;
    END
  END Q2[17]
  PIN Q2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 461.04 13 461.7 13.66 ;
      LAYER Metal4 ;
        RECT 461.04 13 461.7 13.66 ;
      LAYER Metal5 ;
        RECT 461.04 13 461.7 13.66 ;
      LAYER Metal6 ;
        RECT 461.04 13 461.7 13.66 ;
    END
  END Q2[18]
  PIN Q2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 479.44 13 480.1 13.66 ;
      LAYER Metal4 ;
        RECT 479.44 13 480.1 13.66 ;
      LAYER Metal5 ;
        RECT 479.44 13 480.1 13.66 ;
      LAYER Metal6 ;
        RECT 479.44 13 480.1 13.66 ;
    END
  END Q2[19]
  PIN Q2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 45.77 13 46.43 13.66 ;
      LAYER Metal4 ;
        RECT 45.77 13 46.43 13.66 ;
      LAYER Metal5 ;
        RECT 45.77 13 46.43 13.66 ;
      LAYER Metal6 ;
        RECT 45.77 13 46.43 13.66 ;
    END
  END Q2[1]
  PIN Q2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 503.6 13 504.26 13.66 ;
      LAYER Metal4 ;
        RECT 503.6 13 504.26 13.66 ;
      LAYER Metal5 ;
        RECT 503.6 13 504.26 13.66 ;
      LAYER Metal6 ;
        RECT 503.6 13 504.26 13.66 ;
    END
  END Q2[20]
  PIN Q2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 522 13 522.66 13.66 ;
      LAYER Metal4 ;
        RECT 522 13 522.66 13.66 ;
      LAYER Metal5 ;
        RECT 522 13 522.66 13.66 ;
      LAYER Metal6 ;
        RECT 522 13 522.66 13.66 ;
    END
  END Q2[21]
  PIN Q2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 546.16 13 546.82 13.66 ;
      LAYER Metal4 ;
        RECT 546.16 13 546.82 13.66 ;
      LAYER Metal5 ;
        RECT 546.16 13 546.82 13.66 ;
      LAYER Metal6 ;
        RECT 546.16 13 546.82 13.66 ;
    END
  END Q2[22]
  PIN Q2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 564.56 13 565.22 13.66 ;
      LAYER Metal4 ;
        RECT 564.56 13 565.22 13.66 ;
      LAYER Metal5 ;
        RECT 564.56 13 565.22 13.66 ;
      LAYER Metal6 ;
        RECT 564.56 13 565.22 13.66 ;
    END
  END Q2[23]
  PIN Q2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 588.72 13 589.38 13.66 ;
      LAYER Metal4 ;
        RECT 588.72 13 589.38 13.66 ;
      LAYER Metal5 ;
        RECT 588.72 13 589.38 13.66 ;
      LAYER Metal6 ;
        RECT 588.72 13 589.38 13.66 ;
    END
  END Q2[24]
  PIN Q2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 607.12 13 607.78 13.66 ;
      LAYER Metal4 ;
        RECT 607.12 13 607.78 13.66 ;
      LAYER Metal5 ;
        RECT 607.12 13 607.78 13.66 ;
      LAYER Metal6 ;
        RECT 607.12 13 607.78 13.66 ;
    END
  END Q2[25]
  PIN Q2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 631.28 13 631.94 13.66 ;
      LAYER Metal4 ;
        RECT 631.28 13 631.94 13.66 ;
      LAYER Metal5 ;
        RECT 631.28 13 631.94 13.66 ;
      LAYER Metal6 ;
        RECT 631.28 13 631.94 13.66 ;
    END
  END Q2[26]
  PIN Q2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 649.68 13 650.34 13.66 ;
      LAYER Metal4 ;
        RECT 649.68 13 650.34 13.66 ;
      LAYER Metal5 ;
        RECT 649.68 13 650.34 13.66 ;
      LAYER Metal6 ;
        RECT 649.68 13 650.34 13.66 ;
    END
  END Q2[27]
  PIN Q2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 673.84 13 674.5 13.66 ;
      LAYER Metal4 ;
        RECT 673.84 13 674.5 13.66 ;
      LAYER Metal5 ;
        RECT 673.84 13 674.5 13.66 ;
      LAYER Metal6 ;
        RECT 673.84 13 674.5 13.66 ;
    END
  END Q2[28]
  PIN Q2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 692.24 13 692.9 13.66 ;
      LAYER Metal4 ;
        RECT 692.24 13 692.9 13.66 ;
      LAYER Metal5 ;
        RECT 692.24 13 692.9 13.66 ;
      LAYER Metal6 ;
        RECT 692.24 13 692.9 13.66 ;
    END
  END Q2[29]
  PIN Q2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 69.93 13 70.59 13.66 ;
      LAYER Metal4 ;
        RECT 69.93 13 70.59 13.66 ;
      LAYER Metal5 ;
        RECT 69.93 13 70.59 13.66 ;
      LAYER Metal6 ;
        RECT 69.93 13 70.59 13.66 ;
    END
  END Q2[2]
  PIN Q2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 716.4 13 717.06 13.66 ;
      LAYER Metal4 ;
        RECT 716.4 13 717.06 13.66 ;
      LAYER Metal5 ;
        RECT 716.4 13 717.06 13.66 ;
      LAYER Metal6 ;
        RECT 716.4 13 717.06 13.66 ;
    END
  END Q2[30]
  PIN Q2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 734.8 13 735.46 13.66 ;
      LAYER Metal4 ;
        RECT 734.8 13 735.46 13.66 ;
      LAYER Metal5 ;
        RECT 734.8 13 735.46 13.66 ;
      LAYER Metal6 ;
        RECT 734.8 13 735.46 13.66 ;
    END
  END Q2[31]
  PIN Q2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 88.33 13 88.99 13.66 ;
      LAYER Metal4 ;
        RECT 88.33 13 88.99 13.66 ;
      LAYER Metal5 ;
        RECT 88.33 13 88.99 13.66 ;
      LAYER Metal6 ;
        RECT 88.33 13 88.99 13.66 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 112.49 13 113.15 13.66 ;
      LAYER Metal4 ;
        RECT 112.49 13 113.15 13.66 ;
      LAYER Metal5 ;
        RECT 112.49 13 113.15 13.66 ;
      LAYER Metal6 ;
        RECT 112.49 13 113.15 13.66 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 130.89 13 131.55 13.66 ;
      LAYER Metal4 ;
        RECT 130.89 13 131.55 13.66 ;
      LAYER Metal5 ;
        RECT 130.89 13 131.55 13.66 ;
      LAYER Metal6 ;
        RECT 130.89 13 131.55 13.66 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 155.05 13 155.71 13.66 ;
      LAYER Metal4 ;
        RECT 155.05 13 155.71 13.66 ;
      LAYER Metal5 ;
        RECT 155.05 13 155.71 13.66 ;
      LAYER Metal6 ;
        RECT 155.05 13 155.71 13.66 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 173.45 13 174.11 13.66 ;
      LAYER Metal4 ;
        RECT 173.45 13 174.11 13.66 ;
      LAYER Metal5 ;
        RECT 173.45 13 174.11 13.66 ;
      LAYER Metal6 ;
        RECT 173.45 13 174.11 13.66 ;
    END
  END Q2[7]
  PIN Q2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 197.61 13 198.27 13.66 ;
      LAYER Metal4 ;
        RECT 197.61 13 198.27 13.66 ;
      LAYER Metal5 ;
        RECT 197.61 13 198.27 13.66 ;
      LAYER Metal6 ;
        RECT 197.61 13 198.27 13.66 ;
    END
  END Q2[8]
  PIN Q2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 216.01 13 216.67 13.66 ;
      LAYER Metal4 ;
        RECT 216.01 13 216.67 13.66 ;
      LAYER Metal5 ;
        RECT 216.01 13 216.67 13.66 ;
      LAYER Metal6 ;
        RECT 216.01 13 216.67 13.66 ;
    END
  END Q2[9]
  PIN WE1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 397.97 13 398.63 13.66 ;
      LAYER Metal4 ;
        RECT 397.97 13 398.63 13.66 ;
      LAYER Metal5 ;
        RECT 397.97 13 398.63 13.66 ;
      LAYER Metal6 ;
        RECT 397.97 13 398.63 13.66 ;
    END
  END WE1
  PIN WE2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 364.2 13 364.86 13.66 ;
      LAYER Metal4 ;
        RECT 364.2 13 364.86 13.66 ;
      LAYER Metal5 ;
        RECT 364.2 13 364.86 13.66 ;
      LAYER Metal6 ;
        RECT 364.2 13 364.86 13.66 ;
    END
  END WE2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 942.445 806.03 947.445 ;
        RECT 0 0 806.03 5 ;
      LAYER Metal2 ;
        RECT 801.03 0 806.03 947.445 ;
        RECT 0 0 5 947.445 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 936.845 800.43 941.845 ;
        RECT 5.6 5.6 800.43 10.6 ;
      LAYER Metal2 ;
        RECT 795.43 5.6 800.43 941.845 ;
        RECT 5.6 5.6 10.6 941.845 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12.8 13 793.2 935.02 ;
    LAYER Metal2 ;
      RECT 12.8 13 793.2 935.02 ;
    LAYER Metal3 ;
      RECT 12.8 13 793.2 935.02 ;
    LAYER Metal4 ;
      RECT 12.8 13 793.2 935.02 ;
    LAYER Metal5 ;
      RECT 12.8 13 793.2 935.02 ;
    LAYER Metal6 ;
      RECT 12.8 13 793.2 935.02 ;
  END
END MEM2_4096X32

END LIBRARY
