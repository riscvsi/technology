VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO MEM1_1024X32
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN MEM1_1024X32 0 0 ;
  SIZE 436.145 BY 168.5 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 86.31 12.66 86.97 ;
      LAYER Metal6 ;
        RECT 12 86.31 12.66 86.97 ;
      LAYER Metal3 ;
        RECT 12 86.31 12.66 86.97 ;
      LAYER Metal4 ;
        RECT 12 86.31 12.66 86.97 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 80.19 12.66 80.85 ;
      LAYER Metal6 ;
        RECT 12 80.19 12.66 80.85 ;
      LAYER Metal3 ;
        RECT 12 80.19 12.66 80.85 ;
      LAYER Metal4 ;
        RECT 12 80.19 12.66 80.85 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 77.09 12.66 77.75 ;
      LAYER Metal6 ;
        RECT 12 77.09 12.66 77.75 ;
      LAYER Metal3 ;
        RECT 12 77.09 12.66 77.75 ;
      LAYER Metal4 ;
        RECT 12 77.09 12.66 77.75 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 70.97 12.66 71.63 ;
      LAYER Metal6 ;
        RECT 12 70.97 12.66 71.63 ;
      LAYER Metal3 ;
        RECT 12 70.97 12.66 71.63 ;
      LAYER Metal4 ;
        RECT 12 70.97 12.66 71.63 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 67.95 12.66 68.61 ;
      LAYER Metal6 ;
        RECT 12 67.95 12.66 68.61 ;
      LAYER Metal3 ;
        RECT 12 67.95 12.66 68.61 ;
      LAYER Metal4 ;
        RECT 12 67.95 12.66 68.61 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 64.85 12.66 65.51 ;
      LAYER Metal6 ;
        RECT 12 64.85 12.66 65.51 ;
      LAYER Metal3 ;
        RECT 12 64.85 12.66 65.51 ;
      LAYER Metal4 ;
        RECT 12 64.85 12.66 65.51 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 58.73 12.66 59.39 ;
      LAYER Metal6 ;
        RECT 12 58.73 12.66 59.39 ;
      LAYER Metal3 ;
        RECT 12 58.73 12.66 59.39 ;
      LAYER Metal4 ;
        RECT 12 58.73 12.66 59.39 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 55.71 12.66 56.37 ;
      LAYER Metal6 ;
        RECT 12 55.71 12.66 56.37 ;
      LAYER Metal3 ;
        RECT 12 55.71 12.66 56.37 ;
      LAYER Metal4 ;
        RECT 12 55.71 12.66 56.37 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 52.61 12.66 53.27 ;
      LAYER Metal6 ;
        RECT 12 52.61 12.66 53.27 ;
      LAYER Metal3 ;
        RECT 12 52.61 12.66 53.27 ;
      LAYER Metal4 ;
        RECT 12 52.61 12.66 53.27 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 12 46.49 12.66 47.15 ;
      LAYER Metal6 ;
        RECT 12 46.49 12.66 47.15 ;
      LAYER Metal3 ;
        RECT 12 46.49 12.66 47.15 ;
      LAYER Metal4 ;
        RECT 12 46.49 12.66 47.15 ;
    END
  END A[9]
  PIN CE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 237.615 12 238.275 12.66 ;
      LAYER Metal6 ;
        RECT 237.615 12 238.275 12.66 ;
      LAYER Metal3 ;
        RECT 237.615 12 238.275 12.66 ;
      LAYER Metal4 ;
        RECT 237.615 12 238.275 12.66 ;
    END
  END CE
  PIN CK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER Metal5 ;
        RECT 247.36 12 248.02 12.66 ;
      LAYER Metal6 ;
        RECT 247.36 12 248.02 12.66 ;
      LAYER Metal3 ;
        RECT 247.36 12 248.02 12.66 ;
      LAYER Metal4 ;
        RECT 247.36 12 248.02 12.66 ;
    END
  END CK
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 20.48 12 21.14 12.66 ;
      LAYER Metal6 ;
        RECT 20.48 12 21.14 12.66 ;
      LAYER Metal3 ;
        RECT 20.48 12 21.14 12.66 ;
      LAYER Metal4 ;
        RECT 20.48 12 21.14 12.66 ;
    END
  END D[0]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 129 12 129.66 12.66 ;
      LAYER Metal6 ;
        RECT 129 12 129.66 12.66 ;
      LAYER Metal3 ;
        RECT 129 12 129.66 12.66 ;
      LAYER Metal4 ;
        RECT 129 12 129.66 12.66 ;
    END
  END D[10]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 137.04 12 137.7 12.66 ;
      LAYER Metal6 ;
        RECT 137.04 12 137.7 12.66 ;
      LAYER Metal3 ;
        RECT 137.04 12 137.7 12.66 ;
      LAYER Metal4 ;
        RECT 137.04 12 137.7 12.66 ;
    END
  END D[11]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 151.34 12 152 12.66 ;
      LAYER Metal6 ;
        RECT 151.34 12 152 12.66 ;
      LAYER Metal3 ;
        RECT 151.34 12 152 12.66 ;
      LAYER Metal4 ;
        RECT 151.34 12 152 12.66 ;
    END
  END D[12]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 159.38 12 160.04 12.66 ;
      LAYER Metal6 ;
        RECT 159.38 12 160.04 12.66 ;
      LAYER Metal3 ;
        RECT 159.38 12 160.04 12.66 ;
      LAYER Metal4 ;
        RECT 159.38 12 160.04 12.66 ;
    END
  END D[13]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 172.62 12 173.28 12.66 ;
      LAYER Metal6 ;
        RECT 172.62 12 173.28 12.66 ;
      LAYER Metal3 ;
        RECT 172.62 12 173.28 12.66 ;
      LAYER Metal4 ;
        RECT 172.62 12 173.28 12.66 ;
    END
  END D[14]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 180.66 12 181.32 12.66 ;
      LAYER Metal6 ;
        RECT 180.66 12 181.32 12.66 ;
      LAYER Metal3 ;
        RECT 180.66 12 181.32 12.66 ;
      LAYER Metal4 ;
        RECT 180.66 12 181.32 12.66 ;
    END
  END D[15]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 254.825 12 255.485 12.66 ;
      LAYER Metal6 ;
        RECT 254.825 12 255.485 12.66 ;
      LAYER Metal3 ;
        RECT 254.825 12 255.485 12.66 ;
      LAYER Metal4 ;
        RECT 254.825 12 255.485 12.66 ;
    END
  END D[16]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 262.865 12 263.525 12.66 ;
      LAYER Metal6 ;
        RECT 262.865 12 263.525 12.66 ;
      LAYER Metal3 ;
        RECT 262.865 12 263.525 12.66 ;
      LAYER Metal4 ;
        RECT 262.865 12 263.525 12.66 ;
    END
  END D[17]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 276.105 12 276.765 12.66 ;
      LAYER Metal6 ;
        RECT 276.105 12 276.765 12.66 ;
      LAYER Metal3 ;
        RECT 276.105 12 276.765 12.66 ;
      LAYER Metal4 ;
        RECT 276.105 12 276.765 12.66 ;
    END
  END D[18]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 284.145 12 284.805 12.66 ;
      LAYER Metal6 ;
        RECT 284.145 12 284.805 12.66 ;
      LAYER Metal3 ;
        RECT 284.145 12 284.805 12.66 ;
      LAYER Metal4 ;
        RECT 284.145 12 284.805 12.66 ;
    END
  END D[19]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 28.52 12 29.18 12.66 ;
      LAYER Metal6 ;
        RECT 28.52 12 29.18 12.66 ;
      LAYER Metal3 ;
        RECT 28.52 12 29.18 12.66 ;
      LAYER Metal4 ;
        RECT 28.52 12 29.18 12.66 ;
    END
  END D[1]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 298.445 12 299.105 12.66 ;
      LAYER Metal6 ;
        RECT 298.445 12 299.105 12.66 ;
      LAYER Metal3 ;
        RECT 298.445 12 299.105 12.66 ;
      LAYER Metal4 ;
        RECT 298.445 12 299.105 12.66 ;
    END
  END D[20]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 306.485 12 307.145 12.66 ;
      LAYER Metal6 ;
        RECT 306.485 12 307.145 12.66 ;
      LAYER Metal3 ;
        RECT 306.485 12 307.145 12.66 ;
      LAYER Metal4 ;
        RECT 306.485 12 307.145 12.66 ;
    END
  END D[21]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 319.725 12 320.385 12.66 ;
      LAYER Metal6 ;
        RECT 319.725 12 320.385 12.66 ;
      LAYER Metal3 ;
        RECT 319.725 12 320.385 12.66 ;
      LAYER Metal4 ;
        RECT 319.725 12 320.385 12.66 ;
    END
  END D[22]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 327.765 12 328.425 12.66 ;
      LAYER Metal6 ;
        RECT 327.765 12 328.425 12.66 ;
      LAYER Metal3 ;
        RECT 327.765 12 328.425 12.66 ;
      LAYER Metal4 ;
        RECT 327.765 12 328.425 12.66 ;
    END
  END D[23]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 342.065 12 342.725 12.66 ;
      LAYER Metal6 ;
        RECT 342.065 12 342.725 12.66 ;
      LAYER Metal3 ;
        RECT 342.065 12 342.725 12.66 ;
      LAYER Metal4 ;
        RECT 342.065 12 342.725 12.66 ;
    END
  END D[24]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 350.105 12 350.765 12.66 ;
      LAYER Metal6 ;
        RECT 350.105 12 350.765 12.66 ;
      LAYER Metal3 ;
        RECT 350.105 12 350.765 12.66 ;
      LAYER Metal4 ;
        RECT 350.105 12 350.765 12.66 ;
    END
  END D[25]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 363.345 12 364.005 12.66 ;
      LAYER Metal6 ;
        RECT 363.345 12 364.005 12.66 ;
      LAYER Metal3 ;
        RECT 363.345 12 364.005 12.66 ;
      LAYER Metal4 ;
        RECT 363.345 12 364.005 12.66 ;
    END
  END D[26]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 371.385 12 372.045 12.66 ;
      LAYER Metal6 ;
        RECT 371.385 12 372.045 12.66 ;
      LAYER Metal3 ;
        RECT 371.385 12 372.045 12.66 ;
      LAYER Metal4 ;
        RECT 371.385 12 372.045 12.66 ;
    END
  END D[27]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 385.685 12 386.345 12.66 ;
      LAYER Metal6 ;
        RECT 385.685 12 386.345 12.66 ;
      LAYER Metal3 ;
        RECT 385.685 12 386.345 12.66 ;
      LAYER Metal4 ;
        RECT 385.685 12 386.345 12.66 ;
    END
  END D[28]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 393.725 12 394.385 12.66 ;
      LAYER Metal6 ;
        RECT 393.725 12 394.385 12.66 ;
      LAYER Metal3 ;
        RECT 393.725 12 394.385 12.66 ;
      LAYER Metal4 ;
        RECT 393.725 12 394.385 12.66 ;
    END
  END D[29]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 41.76 12 42.42 12.66 ;
      LAYER Metal6 ;
        RECT 41.76 12 42.42 12.66 ;
      LAYER Metal3 ;
        RECT 41.76 12 42.42 12.66 ;
      LAYER Metal4 ;
        RECT 41.76 12 42.42 12.66 ;
    END
  END D[2]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 406.965 12 407.625 12.66 ;
      LAYER Metal6 ;
        RECT 406.965 12 407.625 12.66 ;
      LAYER Metal3 ;
        RECT 406.965 12 407.625 12.66 ;
      LAYER Metal4 ;
        RECT 406.965 12 407.625 12.66 ;
    END
  END D[30]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 415.005 12 415.665 12.66 ;
      LAYER Metal6 ;
        RECT 415.005 12 415.665 12.66 ;
      LAYER Metal3 ;
        RECT 415.005 12 415.665 12.66 ;
      LAYER Metal4 ;
        RECT 415.005 12 415.665 12.66 ;
    END
  END D[31]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 49.8 12 50.46 12.66 ;
      LAYER Metal6 ;
        RECT 49.8 12 50.46 12.66 ;
      LAYER Metal3 ;
        RECT 49.8 12 50.46 12.66 ;
      LAYER Metal4 ;
        RECT 49.8 12 50.46 12.66 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 64.1 12 64.76 12.66 ;
      LAYER Metal6 ;
        RECT 64.1 12 64.76 12.66 ;
      LAYER Metal3 ;
        RECT 64.1 12 64.76 12.66 ;
      LAYER Metal4 ;
        RECT 64.1 12 64.76 12.66 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 72.14 12 72.8 12.66 ;
      LAYER Metal6 ;
        RECT 72.14 12 72.8 12.66 ;
      LAYER Metal3 ;
        RECT 72.14 12 72.8 12.66 ;
      LAYER Metal4 ;
        RECT 72.14 12 72.8 12.66 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 85.38 12 86.04 12.66 ;
      LAYER Metal6 ;
        RECT 85.38 12 86.04 12.66 ;
      LAYER Metal3 ;
        RECT 85.38 12 86.04 12.66 ;
      LAYER Metal4 ;
        RECT 85.38 12 86.04 12.66 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 93.42 12 94.08 12.66 ;
      LAYER Metal6 ;
        RECT 93.42 12 94.08 12.66 ;
      LAYER Metal3 ;
        RECT 93.42 12 94.08 12.66 ;
      LAYER Metal4 ;
        RECT 93.42 12 94.08 12.66 ;
    END
  END D[7]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 107.72 12 108.38 12.66 ;
      LAYER Metal6 ;
        RECT 107.72 12 108.38 12.66 ;
      LAYER Metal3 ;
        RECT 107.72 12 108.38 12.66 ;
      LAYER Metal4 ;
        RECT 107.72 12 108.38 12.66 ;
    END
  END D[8]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 115.76 12 116.42 12.66 ;
      LAYER Metal6 ;
        RECT 115.76 12 116.42 12.66 ;
      LAYER Metal3 ;
        RECT 115.76 12 116.42 12.66 ;
      LAYER Metal4 ;
        RECT 115.76 12 116.42 12.66 ;
    END
  END D[9]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 23.06 12 23.72 12.66 ;
      LAYER Metal6 ;
        RECT 23.06 12 23.72 12.66 ;
      LAYER Metal3 ;
        RECT 23.06 12 23.72 12.66 ;
      LAYER Metal4 ;
        RECT 23.06 12 23.72 12.66 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 131.58 12 132.24 12.66 ;
      LAYER Metal6 ;
        RECT 131.58 12 132.24 12.66 ;
      LAYER Metal3 ;
        RECT 131.58 12 132.24 12.66 ;
      LAYER Metal4 ;
        RECT 131.58 12 132.24 12.66 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 134.46 12 135.12 12.66 ;
      LAYER Metal6 ;
        RECT 134.46 12 135.12 12.66 ;
      LAYER Metal3 ;
        RECT 134.46 12 135.12 12.66 ;
      LAYER Metal4 ;
        RECT 134.46 12 135.12 12.66 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 153.92 12 154.58 12.66 ;
      LAYER Metal6 ;
        RECT 153.92 12 154.58 12.66 ;
      LAYER Metal3 ;
        RECT 153.92 12 154.58 12.66 ;
      LAYER Metal4 ;
        RECT 153.92 12 154.58 12.66 ;
    END
  END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 156.8 12 157.46 12.66 ;
      LAYER Metal6 ;
        RECT 156.8 12 157.46 12.66 ;
      LAYER Metal3 ;
        RECT 156.8 12 157.46 12.66 ;
      LAYER Metal4 ;
        RECT 156.8 12 157.46 12.66 ;
    END
  END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 175.2 12 175.86 12.66 ;
      LAYER Metal6 ;
        RECT 175.2 12 175.86 12.66 ;
      LAYER Metal3 ;
        RECT 175.2 12 175.86 12.66 ;
      LAYER Metal4 ;
        RECT 175.2 12 175.86 12.66 ;
    END
  END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 178.08 12 178.74 12.66 ;
      LAYER Metal6 ;
        RECT 178.08 12 178.74 12.66 ;
      LAYER Metal3 ;
        RECT 178.08 12 178.74 12.66 ;
      LAYER Metal4 ;
        RECT 178.08 12 178.74 12.66 ;
    END
  END Q[15]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 257.405 12 258.065 12.66 ;
      LAYER Metal6 ;
        RECT 257.405 12 258.065 12.66 ;
      LAYER Metal3 ;
        RECT 257.405 12 258.065 12.66 ;
      LAYER Metal4 ;
        RECT 257.405 12 258.065 12.66 ;
    END
  END Q[16]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 260.285 12 260.945 12.66 ;
      LAYER Metal6 ;
        RECT 260.285 12 260.945 12.66 ;
      LAYER Metal3 ;
        RECT 260.285 12 260.945 12.66 ;
      LAYER Metal4 ;
        RECT 260.285 12 260.945 12.66 ;
    END
  END Q[17]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 278.685 12 279.345 12.66 ;
      LAYER Metal6 ;
        RECT 278.685 12 279.345 12.66 ;
      LAYER Metal3 ;
        RECT 278.685 12 279.345 12.66 ;
      LAYER Metal4 ;
        RECT 278.685 12 279.345 12.66 ;
    END
  END Q[18]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 281.565 12 282.225 12.66 ;
      LAYER Metal6 ;
        RECT 281.565 12 282.225 12.66 ;
      LAYER Metal3 ;
        RECT 281.565 12 282.225 12.66 ;
      LAYER Metal4 ;
        RECT 281.565 12 282.225 12.66 ;
    END
  END Q[19]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 25.94 12 26.6 12.66 ;
      LAYER Metal6 ;
        RECT 25.94 12 26.6 12.66 ;
      LAYER Metal3 ;
        RECT 25.94 12 26.6 12.66 ;
      LAYER Metal4 ;
        RECT 25.94 12 26.6 12.66 ;
    END
  END Q[1]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 301.025 12 301.685 12.66 ;
      LAYER Metal6 ;
        RECT 301.025 12 301.685 12.66 ;
      LAYER Metal3 ;
        RECT 301.025 12 301.685 12.66 ;
      LAYER Metal4 ;
        RECT 301.025 12 301.685 12.66 ;
    END
  END Q[20]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 303.905 12 304.565 12.66 ;
      LAYER Metal6 ;
        RECT 303.905 12 304.565 12.66 ;
      LAYER Metal3 ;
        RECT 303.905 12 304.565 12.66 ;
      LAYER Metal4 ;
        RECT 303.905 12 304.565 12.66 ;
    END
  END Q[21]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 322.305 12 322.965 12.66 ;
      LAYER Metal6 ;
        RECT 322.305 12 322.965 12.66 ;
      LAYER Metal3 ;
        RECT 322.305 12 322.965 12.66 ;
      LAYER Metal4 ;
        RECT 322.305 12 322.965 12.66 ;
    END
  END Q[22]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 325.185 12 325.845 12.66 ;
      LAYER Metal6 ;
        RECT 325.185 12 325.845 12.66 ;
      LAYER Metal3 ;
        RECT 325.185 12 325.845 12.66 ;
      LAYER Metal4 ;
        RECT 325.185 12 325.845 12.66 ;
    END
  END Q[23]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 344.645 12 345.305 12.66 ;
      LAYER Metal6 ;
        RECT 344.645 12 345.305 12.66 ;
      LAYER Metal3 ;
        RECT 344.645 12 345.305 12.66 ;
      LAYER Metal4 ;
        RECT 344.645 12 345.305 12.66 ;
    END
  END Q[24]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 347.525 12 348.185 12.66 ;
      LAYER Metal6 ;
        RECT 347.525 12 348.185 12.66 ;
      LAYER Metal3 ;
        RECT 347.525 12 348.185 12.66 ;
      LAYER Metal4 ;
        RECT 347.525 12 348.185 12.66 ;
    END
  END Q[25]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 365.925 12 366.585 12.66 ;
      LAYER Metal6 ;
        RECT 365.925 12 366.585 12.66 ;
      LAYER Metal3 ;
        RECT 365.925 12 366.585 12.66 ;
      LAYER Metal4 ;
        RECT 365.925 12 366.585 12.66 ;
    END
  END Q[26]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 368.805 12 369.465 12.66 ;
      LAYER Metal6 ;
        RECT 368.805 12 369.465 12.66 ;
      LAYER Metal3 ;
        RECT 368.805 12 369.465 12.66 ;
      LAYER Metal4 ;
        RECT 368.805 12 369.465 12.66 ;
    END
  END Q[27]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 388.265 12 388.925 12.66 ;
      LAYER Metal6 ;
        RECT 388.265 12 388.925 12.66 ;
      LAYER Metal3 ;
        RECT 388.265 12 388.925 12.66 ;
      LAYER Metal4 ;
        RECT 388.265 12 388.925 12.66 ;
    END
  END Q[28]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 391.145 12 391.805 12.66 ;
      LAYER Metal6 ;
        RECT 391.145 12 391.805 12.66 ;
      LAYER Metal3 ;
        RECT 391.145 12 391.805 12.66 ;
      LAYER Metal4 ;
        RECT 391.145 12 391.805 12.66 ;
    END
  END Q[29]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 44.34 12 45 12.66 ;
      LAYER Metal6 ;
        RECT 44.34 12 45 12.66 ;
      LAYER Metal3 ;
        RECT 44.34 12 45 12.66 ;
      LAYER Metal4 ;
        RECT 44.34 12 45 12.66 ;
    END
  END Q[2]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 409.545 12 410.205 12.66 ;
      LAYER Metal6 ;
        RECT 409.545 12 410.205 12.66 ;
      LAYER Metal3 ;
        RECT 409.545 12 410.205 12.66 ;
      LAYER Metal4 ;
        RECT 409.545 12 410.205 12.66 ;
    END
  END Q[30]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 412.425 12 413.085 12.66 ;
      LAYER Metal6 ;
        RECT 412.425 12 413.085 12.66 ;
      LAYER Metal3 ;
        RECT 412.425 12 413.085 12.66 ;
      LAYER Metal4 ;
        RECT 412.425 12 413.085 12.66 ;
    END
  END Q[31]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 47.22 12 47.88 12.66 ;
      LAYER Metal6 ;
        RECT 47.22 12 47.88 12.66 ;
      LAYER Metal3 ;
        RECT 47.22 12 47.88 12.66 ;
      LAYER Metal4 ;
        RECT 47.22 12 47.88 12.66 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 66.68 12 67.34 12.66 ;
      LAYER Metal6 ;
        RECT 66.68 12 67.34 12.66 ;
      LAYER Metal3 ;
        RECT 66.68 12 67.34 12.66 ;
      LAYER Metal4 ;
        RECT 66.68 12 67.34 12.66 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 69.56 12 70.22 12.66 ;
      LAYER Metal6 ;
        RECT 69.56 12 70.22 12.66 ;
      LAYER Metal3 ;
        RECT 69.56 12 70.22 12.66 ;
      LAYER Metal4 ;
        RECT 69.56 12 70.22 12.66 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 87.96 12 88.62 12.66 ;
      LAYER Metal6 ;
        RECT 87.96 12 88.62 12.66 ;
      LAYER Metal3 ;
        RECT 87.96 12 88.62 12.66 ;
      LAYER Metal4 ;
        RECT 87.96 12 88.62 12.66 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 90.84 12 91.5 12.66 ;
      LAYER Metal6 ;
        RECT 90.84 12 91.5 12.66 ;
      LAYER Metal3 ;
        RECT 90.84 12 91.5 12.66 ;
      LAYER Metal4 ;
        RECT 90.84 12 91.5 12.66 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 110.3 12 110.96 12.66 ;
      LAYER Metal6 ;
        RECT 110.3 12 110.96 12.66 ;
      LAYER Metal3 ;
        RECT 110.3 12 110.96 12.66 ;
      LAYER Metal4 ;
        RECT 110.3 12 110.96 12.66 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 113.18 12 113.84 12.66 ;
      LAYER Metal6 ;
        RECT 113.18 12 113.84 12.66 ;
      LAYER Metal3 ;
        RECT 113.18 12 113.84 12.66 ;
      LAYER Metal4 ;
        RECT 113.18 12 113.84 12.66 ;
    END
  END Q[9]
  PIN WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal5 ;
        RECT 243.66 12 244.32 12.66 ;
      LAYER Metal6 ;
        RECT 243.66 12 244.32 12.66 ;
      LAYER Metal3 ;
        RECT 243.66 12 244.32 12.66 ;
      LAYER Metal4 ;
        RECT 243.66 12 244.32 12.66 ;
    END
  END WE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 0 163.5 436.145 168.5 ;
        RECT 0 0 436.145 5 ;
      LAYER Metal2 ;
        RECT 431.145 0 436.145 168.5 ;
        RECT 0 0 5 168.5 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER Metal1 ;
        RECT 5.6 157.9 430.545 162.9 ;
        RECT 5.6 5.6 430.545 10.6 ;
      LAYER Metal2 ;
        RECT 425.545 5.6 430.545 162.9 ;
        RECT 5.6 5.6 10.6 162.9 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 12 12 424.135 156.495 ;
    LAYER Metal2 ;
      RECT 12 12 424.135 156.495 ;
    LAYER Metal3 ;
      RECT 12 12 424.135 156.495 ;
    LAYER Metal4 ;
      RECT 12 12 424.135 156.495 ;
    LAYER Metal5 ;
      RECT 12 12 424.135 156.495 ;
    LAYER Metal6 ;
      RECT 12 12 424.135 156.495 ;
  END
END MEM1_1024X32

END LIBRARY
